magic
tech sky130A
timestamp 1616960036
<< nwell >>
rect 0 324 308 503
rect 66 300 240 324
rect 141 239 240 300
<< nmos >>
rect 47 223 62 265
rect 53 72 68 172
rect 203 156 245 171
rect 203 105 245 120
<< pmos >>
rect 78 346 93 401
rect 165 381 265 396
rect 165 291 220 306
<< ndiff >>
rect 7 253 47 265
rect 7 236 17 253
rect 34 236 47 253
rect 7 223 47 236
rect 62 253 107 265
rect 62 236 77 253
rect 94 236 107 253
rect 62 223 107 236
rect 203 197 245 205
rect 8 161 53 172
rect 8 144 21 161
rect 38 144 53 161
rect 8 118 53 144
rect 8 101 21 118
rect 38 101 53 118
rect 8 72 53 101
rect 68 143 108 172
rect 203 180 215 197
rect 232 180 245 197
rect 203 171 245 180
rect 68 126 82 143
rect 99 126 108 143
rect 68 102 108 126
rect 203 147 245 156
rect 203 130 215 147
rect 232 130 245 147
rect 203 120 245 130
rect 68 85 82 102
rect 99 85 108 102
rect 68 72 108 85
rect 203 95 245 105
rect 203 78 215 95
rect 232 78 245 95
rect 203 70 245 78
<< pdiff >>
rect 165 423 265 433
rect 165 406 202 423
rect 219 406 237 423
rect 254 406 265 423
rect 38 382 78 401
rect 38 365 48 382
rect 65 365 78 382
rect 38 346 78 365
rect 93 382 138 401
rect 165 396 265 406
rect 93 365 108 382
rect 125 365 138 382
rect 93 346 138 365
rect 165 372 265 381
rect 165 355 184 372
rect 201 355 237 372
rect 254 355 265 372
rect 165 342 265 355
rect 165 332 220 342
rect 165 315 184 332
rect 201 315 220 332
rect 165 306 220 315
rect 165 282 220 291
rect 165 265 184 282
rect 201 265 220 282
rect 165 257 220 265
<< ndiffc >>
rect 17 236 34 253
rect 77 236 94 253
rect 21 144 38 161
rect 21 101 38 118
rect 215 180 232 197
rect 82 126 99 143
rect 215 130 232 147
rect 82 85 99 102
rect 215 78 232 95
<< pdiffc >>
rect 202 406 219 423
rect 237 406 254 423
rect 48 365 65 382
rect 108 365 125 382
rect 184 355 201 372
rect 237 355 254 372
rect 184 315 201 332
rect 184 265 201 282
<< psubdiff >>
rect 38 8 79 20
rect 38 -9 50 8
rect 67 -9 79 8
rect 38 -21 79 -9
<< nsubdiff >>
rect 19 467 72 485
rect 19 450 37 467
rect 54 450 72 467
rect 19 432 72 450
<< psubdiffcont >>
rect 50 -9 67 8
<< nsubdiffcont >>
rect 37 450 54 467
<< poly >>
rect 78 401 93 418
rect 152 381 165 396
rect 265 381 295 396
rect 78 329 93 346
rect 78 321 117 329
rect 78 304 92 321
rect 109 304 117 321
rect 280 306 295 381
rect 78 296 117 304
rect 78 294 93 296
rect 47 279 93 294
rect 152 291 165 306
rect 220 298 295 306
rect 220 291 270 298
rect 47 265 62 279
rect 262 281 270 291
rect 287 281 295 298
rect 262 273 295 281
rect 47 208 62 223
rect 260 222 293 230
rect 260 205 268 222
rect 285 205 293 222
rect 260 197 293 205
rect 53 172 68 186
rect 126 181 159 189
rect 126 164 134 181
rect 151 171 159 181
rect 151 164 203 171
rect 126 156 203 164
rect 245 156 260 171
rect 135 155 150 156
rect 258 121 291 129
rect 258 120 266 121
rect 180 105 203 120
rect 245 105 266 120
rect 258 104 266 105
rect 283 104 291 121
rect 258 96 291 104
rect 53 58 68 72
rect 126 58 159 66
rect 53 43 134 58
rect 126 41 134 43
rect 151 41 159 58
rect 126 33 159 41
<< polycont >>
rect 92 304 109 321
rect 270 281 287 298
rect 268 205 285 222
rect 134 164 151 181
rect 266 104 283 121
rect 134 41 151 58
<< locali >>
rect 29 467 62 475
rect 0 450 37 467
rect 54 450 308 467
rect 29 442 62 450
rect 100 390 117 450
rect 176 423 262 431
rect 176 406 202 423
rect 219 406 237 423
rect 254 406 262 423
rect 176 398 262 406
rect 40 382 73 390
rect 40 365 48 382
rect 65 365 73 382
rect 40 357 73 365
rect 100 382 133 390
rect 100 365 108 382
rect 125 365 133 382
rect 100 357 133 365
rect 176 372 262 380
rect 48 328 65 357
rect 176 355 184 372
rect 201 355 237 372
rect 254 355 262 372
rect 176 347 262 355
rect 176 332 209 347
rect 25 311 65 328
rect 84 321 136 329
rect 25 294 42 311
rect 84 304 92 321
rect 109 304 136 321
rect 176 315 184 332
rect 201 315 209 332
rect 176 307 209 315
rect 84 296 136 304
rect 14 288 42 294
rect 14 271 20 288
rect 37 271 42 288
rect 14 265 42 271
rect 9 253 42 265
rect 9 236 17 253
rect 34 236 42 253
rect 9 228 42 236
rect 69 253 102 261
rect 69 236 77 253
rect 94 236 102 253
rect 69 228 102 236
rect 119 234 136 296
rect 262 298 295 306
rect 176 282 209 290
rect 176 265 184 282
rect 201 277 209 282
rect 262 281 270 298
rect 287 281 295 298
rect 262 277 295 281
rect 201 265 295 277
rect 176 257 295 265
rect 215 239 232 257
rect 13 161 46 169
rect 13 144 21 161
rect 38 144 46 161
rect 80 154 100 228
rect 119 217 196 234
rect 260 222 293 230
rect 179 205 196 217
rect 260 205 268 222
rect 285 205 293 222
rect 179 197 240 205
rect 260 197 293 205
rect 126 181 159 189
rect 179 182 215 197
rect 126 164 134 181
rect 151 164 159 181
rect 210 180 215 182
rect 232 180 240 197
rect 210 172 240 180
rect 126 156 159 164
rect 13 118 46 144
rect 13 101 21 118
rect 38 101 46 118
rect 13 93 46 101
rect 74 143 107 154
rect 207 147 240 155
rect 74 126 82 143
rect 99 126 107 143
rect 197 130 215 147
rect 232 130 240 147
rect 74 102 107 126
rect 207 122 240 130
rect 268 129 285 197
rect 258 121 291 129
rect 258 104 266 121
rect 283 104 291 121
rect 74 85 82 102
rect 99 85 107 102
rect 74 77 107 85
rect 90 8 107 77
rect 207 95 240 103
rect 258 96 291 104
rect 207 78 215 95
rect 232 78 240 95
rect 207 70 240 78
rect 126 58 159 66
rect 126 41 134 58
rect 151 41 159 58
rect 126 33 159 41
rect 0 -9 50 8
rect 67 -9 308 8
<< viali >>
rect 37 450 54 467
rect 202 406 219 423
rect 237 355 254 372
rect 92 304 109 321
rect 20 271 37 288
rect 21 144 38 161
rect 215 222 232 239
rect 268 205 285 222
rect 134 164 151 181
rect 21 101 38 118
rect 180 130 197 147
rect 215 78 232 95
rect 134 41 151 58
rect 50 -9 67 8
<< metal1 >>
rect 0 444 31 473
rect 60 444 308 473
rect 196 423 225 429
rect 196 406 202 423
rect 219 406 225 423
rect 196 400 225 406
rect 196 347 210 400
rect 240 378 260 444
rect 231 372 260 378
rect 231 355 237 372
rect 254 355 260 372
rect 231 349 260 355
rect 101 329 210 347
rect 100 327 117 329
rect 86 321 117 327
rect 86 304 92 321
rect 109 320 117 321
rect 109 304 115 320
rect 86 298 115 304
rect 14 288 42 294
rect 14 284 20 288
rect 0 271 20 284
rect 37 284 42 288
rect 37 271 308 284
rect 0 267 308 271
rect 14 265 42 267
rect 209 239 238 245
rect 209 222 215 239
rect 232 222 238 239
rect 209 216 238 222
rect 259 228 294 231
rect 125 187 160 190
rect 15 161 46 167
rect 15 144 21 161
rect 38 144 46 161
rect 125 158 128 187
rect 157 158 160 187
rect 125 155 160 158
rect 15 138 46 144
rect 174 147 203 153
rect 174 138 180 147
rect 15 130 180 138
rect 197 130 203 147
rect 15 124 203 130
rect 15 118 46 124
rect 15 101 21 118
rect 38 101 46 118
rect 220 101 235 216
rect 259 199 262 228
rect 291 199 294 228
rect 259 196 294 199
rect 15 95 46 101
rect 209 95 238 101
rect 209 78 215 95
rect 232 78 238 95
rect 209 72 238 78
rect 128 58 157 64
rect 0 41 134 58
rect 151 41 308 58
rect 126 33 159 41
rect 0 -15 43 14
rect 72 -15 308 14
<< via1 >>
rect 31 467 60 473
rect 31 450 37 467
rect 37 450 54 467
rect 54 450 60 467
rect 31 444 60 450
rect 128 181 157 187
rect 128 164 134 181
rect 134 164 151 181
rect 151 164 157 181
rect 128 158 157 164
rect 262 222 291 228
rect 262 205 268 222
rect 268 205 285 222
rect 285 205 291 222
rect 262 199 291 205
rect 43 8 72 14
rect 43 -9 50 8
rect 50 -9 67 8
rect 67 -9 72 8
rect 43 -15 72 -9
<< metal2 >>
rect 23 476 68 481
rect 23 441 28 476
rect 63 441 68 476
rect 23 436 68 441
rect 134 190 151 503
rect 268 231 285 503
rect 259 228 294 231
rect 259 199 262 228
rect 291 199 294 228
rect 259 196 294 199
rect 125 187 160 190
rect 125 158 128 187
rect 157 158 160 187
rect 125 155 160 158
rect 35 17 80 22
rect 35 -18 40 17
rect 75 -18 80 17
rect 35 -23 80 -18
rect 134 -25 151 155
rect 268 -25 285 196
<< via2 >>
rect 28 473 63 476
rect 28 444 31 473
rect 31 444 60 473
rect 60 444 63 473
rect 28 441 63 444
rect 40 14 75 17
rect 40 -15 43 14
rect 43 -15 72 14
rect 72 -15 75 14
rect 40 -18 75 -15
<< metal3 >>
rect 19 476 72 485
rect 0 441 28 476
rect 63 441 308 476
rect 19 432 72 441
rect 30 17 82 25
rect 30 15 40 17
rect 0 -15 40 15
rect 30 -18 40 -15
rect 75 15 82 17
rect 75 -15 308 15
rect 75 -18 82 -15
rect 30 -25 82 -18
<< labels >>
flabel metal2 s 130 161 154 185 0 FreeSans 200 0 0 0 bl
port 0 nsew
flabel metal2 s 264 202 288 226 0 FreeSans 200 0 0 0 br
port 1 nsew
flabel metal1 s 17 269 41 293 0 FreeSans 200 0 0 0 dout
port 2 nsew
flabel metal3 s 33 447 57 471 0 FreeSans 200 0 0 0 vdd
port 4 nsew
flabel metal3 s 45 -11 69 13 0 FreeSans 200 0 0 0 gnd
port 5 nsew
flabel metal1 s 129 39 153 63 0 FreeSans 200 0 0 0 en
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 308 459
<< end >>
