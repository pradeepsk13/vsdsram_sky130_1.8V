VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_sky130A
   CLASS BLOCK ;
   SIZE 60.17 BY 118.34 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  12.86 -10.1 13.38 -9.58 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  25.16 -10.1 25.68 -9.58 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -11.74 117.82 -11.22 118.34 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -14.2 117.82 -13.68 118.34 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -13.38 117.82 -12.86 118.34 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -12.56 117.82 -12.04 118.34 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  -56.84 -7.64 -56.32 -7.12 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  -56.84 -4.36 -56.32 -3.84 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -24.86 -10.1 -24.34 -9.58 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  59.6 10.4 60.12 10.92 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  59.6 11.22 60.12 11.74 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -56.02 -6.0 -54.68 -4.66 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -56.02 -10.1 -54.68 -8.76 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  52.29 35.41 52.58 35.47 ;
      RECT  52.04 33.58 52.33 33.64 ;
      RECT  49.61 33.64 52.69 33.79 ;
      RECT  50.06 37.37 50.41 37.72 ;
      RECT  50.81 36.41 52.0 36.58 ;
      RECT  52.3 34.32 52.59 34.38 ;
      RECT  50.17 36.5 50.33 37.06 ;
      RECT  51.76 35.38 52.11 35.47 ;
      RECT  50.97 34.32 51.32 34.41 ;
      RECT  50.97 34.06 51.32 34.15 ;
      RECT  50.59 34.56 51.04 34.7 ;
      RECT  51.77 37.08 52.06 37.37 ;
      RECT  51.76 35.47 52.58 35.64 ;
      RECT  51.03 37.22 51.32 37.37 ;
      RECT  51.83 36.58 52.0 37.08 ;
      RECT  50.87 34.7 51.04 36.35 ;
      RECT  50.06 33.14 50.41 33.49 ;
      RECT  50.17 37.08 51.32 37.22 ;
      RECT  49.76 36.17 50.33 36.5 ;
      RECT  50.97 34.15 52.59 34.32 ;
      RECT  50.59 34.38 50.76 34.56 ;
      RECT  52.3 34.09 52.59 34.15 ;
      RECT  50.53 34.09 50.82 34.38 ;
      RECT  50.81 36.58 51.1 36.64 ;
      RECT  50.81 36.35 51.1 36.41 ;
      RECT  52.04 33.79 52.33 33.87 ;
      RECT  52.29 35.64 52.58 35.7 ;
      RECT  50.17 37.06 51.04 37.08 ;
      RECT  51.76 35.64 52.11 35.73 ;
      RECT  52.29 39.91 52.58 39.85 ;
      RECT  52.04 41.74 52.33 41.68 ;
      RECT  49.61 41.68 52.69 41.53 ;
      RECT  50.06 37.95 50.41 37.6 ;
      RECT  50.81 38.91 52.0 38.74 ;
      RECT  52.3 41.0 52.59 40.94 ;
      RECT  50.17 38.82 50.33 38.26 ;
      RECT  51.76 39.94 52.11 39.85 ;
      RECT  50.97 41.0 51.32 40.91 ;
      RECT  50.97 41.26 51.32 41.17 ;
      RECT  50.59 40.76 51.04 40.62 ;
      RECT  51.77 38.24 52.06 37.95 ;
      RECT  51.76 39.85 52.58 39.68 ;
      RECT  51.03 38.1 51.32 37.95 ;
      RECT  51.83 38.74 52.0 38.24 ;
      RECT  50.87 40.62 51.04 38.97 ;
      RECT  50.06 42.18 50.41 41.83 ;
      RECT  50.17 38.24 51.32 38.1 ;
      RECT  49.76 39.15 50.33 38.82 ;
      RECT  50.97 41.17 52.59 41.0 ;
      RECT  50.59 40.94 50.76 40.76 ;
      RECT  52.3 41.23 52.59 41.17 ;
      RECT  50.53 41.23 50.82 40.94 ;
      RECT  50.81 38.74 51.1 38.68 ;
      RECT  50.81 38.97 51.1 38.91 ;
      RECT  52.04 41.53 52.33 41.45 ;
      RECT  52.29 39.68 52.58 39.62 ;
      RECT  50.17 38.26 51.04 38.24 ;
      RECT  51.76 39.68 52.11 39.59 ;
      RECT  52.29 44.11 52.58 44.17 ;
      RECT  52.04 42.28 52.33 42.34 ;
      RECT  49.61 42.34 52.69 42.49 ;
      RECT  50.06 46.07 50.41 46.42 ;
      RECT  50.81 45.11 52.0 45.28 ;
      RECT  52.3 43.02 52.59 43.08 ;
      RECT  50.17 45.2 50.33 45.76 ;
      RECT  51.76 44.08 52.11 44.17 ;
      RECT  50.97 43.02 51.32 43.11 ;
      RECT  50.97 42.76 51.32 42.85 ;
      RECT  50.59 43.26 51.04 43.4 ;
      RECT  51.77 45.78 52.06 46.07 ;
      RECT  51.76 44.17 52.58 44.34 ;
      RECT  51.03 45.92 51.32 46.07 ;
      RECT  51.83 45.28 52.0 45.78 ;
      RECT  50.87 43.4 51.04 45.05 ;
      RECT  50.06 41.84 50.41 42.19 ;
      RECT  50.17 45.78 51.32 45.92 ;
      RECT  49.76 44.87 50.33 45.2 ;
      RECT  50.97 42.85 52.59 43.02 ;
      RECT  50.59 43.08 50.76 43.26 ;
      RECT  52.3 42.79 52.59 42.85 ;
      RECT  50.53 42.79 50.82 43.08 ;
      RECT  50.81 45.28 51.1 45.34 ;
      RECT  50.81 45.05 51.1 45.11 ;
      RECT  52.04 42.49 52.33 42.57 ;
      RECT  52.29 44.34 52.58 44.4 ;
      RECT  50.17 45.76 51.04 45.78 ;
      RECT  51.76 44.34 52.11 44.43 ;
      RECT  52.29 48.61 52.58 48.55 ;
      RECT  52.04 50.44 52.33 50.38 ;
      RECT  49.61 50.38 52.69 50.23 ;
      RECT  50.06 46.65 50.41 46.3 ;
      RECT  50.81 47.61 52.0 47.44 ;
      RECT  52.3 49.7 52.59 49.64 ;
      RECT  50.17 47.52 50.33 46.96 ;
      RECT  51.76 48.64 52.11 48.55 ;
      RECT  50.97 49.7 51.32 49.61 ;
      RECT  50.97 49.96 51.32 49.87 ;
      RECT  50.59 49.46 51.04 49.32 ;
      RECT  51.77 46.94 52.06 46.65 ;
      RECT  51.76 48.55 52.58 48.38 ;
      RECT  51.03 46.8 51.32 46.65 ;
      RECT  51.83 47.44 52.0 46.94 ;
      RECT  50.87 49.32 51.04 47.67 ;
      RECT  50.06 50.88 50.41 50.53 ;
      RECT  50.17 46.94 51.32 46.8 ;
      RECT  49.76 47.85 50.33 47.52 ;
      RECT  50.97 49.87 52.59 49.7 ;
      RECT  50.59 49.64 50.76 49.46 ;
      RECT  52.3 49.93 52.59 49.87 ;
      RECT  50.53 49.93 50.82 49.64 ;
      RECT  50.81 47.44 51.1 47.38 ;
      RECT  50.81 47.67 51.1 47.61 ;
      RECT  52.04 50.23 52.33 50.15 ;
      RECT  52.29 48.38 52.58 48.32 ;
      RECT  50.17 46.96 51.04 46.94 ;
      RECT  51.76 48.38 52.11 48.29 ;
      RECT  52.29 52.81 52.58 52.87 ;
      RECT  52.04 50.98 52.33 51.04 ;
      RECT  49.61 51.04 52.69 51.19 ;
      RECT  50.06 54.77 50.41 55.12 ;
      RECT  50.81 53.81 52.0 53.98 ;
      RECT  52.3 51.72 52.59 51.78 ;
      RECT  50.17 53.9 50.33 54.46 ;
      RECT  51.76 52.78 52.11 52.87 ;
      RECT  50.97 51.72 51.32 51.81 ;
      RECT  50.97 51.46 51.32 51.55 ;
      RECT  50.59 51.96 51.04 52.1 ;
      RECT  51.77 54.48 52.06 54.77 ;
      RECT  51.76 52.87 52.58 53.04 ;
      RECT  51.03 54.62 51.32 54.77 ;
      RECT  51.83 53.98 52.0 54.48 ;
      RECT  50.87 52.1 51.04 53.75 ;
      RECT  50.06 50.54 50.41 50.89 ;
      RECT  50.17 54.48 51.32 54.62 ;
      RECT  49.76 53.57 50.33 53.9 ;
      RECT  50.97 51.55 52.59 51.72 ;
      RECT  50.59 51.78 50.76 51.96 ;
      RECT  52.3 51.49 52.59 51.55 ;
      RECT  50.53 51.49 50.82 51.78 ;
      RECT  50.81 53.98 51.1 54.04 ;
      RECT  50.81 53.75 51.1 53.81 ;
      RECT  52.04 51.19 52.33 51.27 ;
      RECT  52.29 53.04 52.58 53.1 ;
      RECT  50.17 54.46 51.04 54.48 ;
      RECT  51.76 53.04 52.11 53.13 ;
      RECT  52.29 57.31 52.58 57.25 ;
      RECT  52.04 59.14 52.33 59.08 ;
      RECT  49.61 59.08 52.69 58.93 ;
      RECT  50.06 55.35 50.41 55.0 ;
      RECT  50.81 56.31 52.0 56.14 ;
      RECT  52.3 58.4 52.59 58.34 ;
      RECT  50.17 56.22 50.33 55.66 ;
      RECT  51.76 57.34 52.11 57.25 ;
      RECT  50.97 58.4 51.32 58.31 ;
      RECT  50.97 58.66 51.32 58.57 ;
      RECT  50.59 58.16 51.04 58.02 ;
      RECT  51.77 55.64 52.06 55.35 ;
      RECT  51.76 57.25 52.58 57.08 ;
      RECT  51.03 55.5 51.32 55.35 ;
      RECT  51.83 56.14 52.0 55.64 ;
      RECT  50.87 58.02 51.04 56.37 ;
      RECT  50.06 59.58 50.41 59.23 ;
      RECT  50.17 55.64 51.32 55.5 ;
      RECT  49.76 56.55 50.33 56.22 ;
      RECT  50.97 58.57 52.59 58.4 ;
      RECT  50.59 58.34 50.76 58.16 ;
      RECT  52.3 58.63 52.59 58.57 ;
      RECT  50.53 58.63 50.82 58.34 ;
      RECT  50.81 56.14 51.1 56.08 ;
      RECT  50.81 56.37 51.1 56.31 ;
      RECT  52.04 58.93 52.33 58.85 ;
      RECT  52.29 57.08 52.58 57.02 ;
      RECT  50.17 55.66 51.04 55.64 ;
      RECT  51.76 57.08 52.11 56.99 ;
      RECT  52.29 61.51 52.58 61.57 ;
      RECT  52.04 59.68 52.33 59.74 ;
      RECT  49.61 59.74 52.69 59.89 ;
      RECT  50.06 63.47 50.41 63.82 ;
      RECT  50.81 62.51 52.0 62.68 ;
      RECT  52.3 60.42 52.59 60.48 ;
      RECT  50.17 62.6 50.33 63.16 ;
      RECT  51.76 61.48 52.11 61.57 ;
      RECT  50.97 60.42 51.32 60.51 ;
      RECT  50.97 60.16 51.32 60.25 ;
      RECT  50.59 60.66 51.04 60.8 ;
      RECT  51.77 63.18 52.06 63.47 ;
      RECT  51.76 61.57 52.58 61.74 ;
      RECT  51.03 63.32 51.32 63.47 ;
      RECT  51.83 62.68 52.0 63.18 ;
      RECT  50.87 60.8 51.04 62.45 ;
      RECT  50.06 59.24 50.41 59.59 ;
      RECT  50.17 63.18 51.32 63.32 ;
      RECT  49.76 62.27 50.33 62.6 ;
      RECT  50.97 60.25 52.59 60.42 ;
      RECT  50.59 60.48 50.76 60.66 ;
      RECT  52.3 60.19 52.59 60.25 ;
      RECT  50.53 60.19 50.82 60.48 ;
      RECT  50.81 62.68 51.1 62.74 ;
      RECT  50.81 62.45 51.1 62.51 ;
      RECT  52.04 59.89 52.33 59.97 ;
      RECT  52.29 61.74 52.58 61.8 ;
      RECT  50.17 63.16 51.04 63.18 ;
      RECT  51.76 61.74 52.11 61.83 ;
      RECT  52.29 66.01 52.58 65.95 ;
      RECT  52.04 67.84 52.33 67.78 ;
      RECT  49.61 67.78 52.69 67.63 ;
      RECT  50.06 64.05 50.41 63.7 ;
      RECT  50.81 65.01 52.0 64.84 ;
      RECT  52.3 67.1 52.59 67.04 ;
      RECT  50.17 64.92 50.33 64.36 ;
      RECT  51.76 66.04 52.11 65.95 ;
      RECT  50.97 67.1 51.32 67.01 ;
      RECT  50.97 67.36 51.32 67.27 ;
      RECT  50.59 66.86 51.04 66.72 ;
      RECT  51.77 64.34 52.06 64.05 ;
      RECT  51.76 65.95 52.58 65.78 ;
      RECT  51.03 64.2 51.32 64.05 ;
      RECT  51.83 64.84 52.0 64.34 ;
      RECT  50.87 66.72 51.04 65.07 ;
      RECT  50.06 68.28 50.41 67.93 ;
      RECT  50.17 64.34 51.32 64.2 ;
      RECT  49.76 65.25 50.33 64.92 ;
      RECT  50.97 67.27 52.59 67.1 ;
      RECT  50.59 67.04 50.76 66.86 ;
      RECT  52.3 67.33 52.59 67.27 ;
      RECT  50.53 67.33 50.82 67.04 ;
      RECT  50.81 64.84 51.1 64.78 ;
      RECT  50.81 65.07 51.1 65.01 ;
      RECT  52.04 67.63 52.33 67.55 ;
      RECT  52.29 65.78 52.58 65.72 ;
      RECT  50.17 64.36 51.04 64.34 ;
      RECT  51.76 65.78 52.11 65.69 ;
      RECT  52.29 70.21 52.58 70.27 ;
      RECT  52.04 68.38 52.33 68.44 ;
      RECT  49.61 68.44 52.69 68.59 ;
      RECT  50.06 72.17 50.41 72.52 ;
      RECT  50.81 71.21 52.0 71.38 ;
      RECT  52.3 69.12 52.59 69.18 ;
      RECT  50.17 71.3 50.33 71.86 ;
      RECT  51.76 70.18 52.11 70.27 ;
      RECT  50.97 69.12 51.32 69.21 ;
      RECT  50.97 68.86 51.32 68.95 ;
      RECT  50.59 69.36 51.04 69.5 ;
      RECT  51.77 71.88 52.06 72.17 ;
      RECT  51.76 70.27 52.58 70.44 ;
      RECT  51.03 72.02 51.32 72.17 ;
      RECT  51.83 71.38 52.0 71.88 ;
      RECT  50.87 69.5 51.04 71.15 ;
      RECT  50.06 67.94 50.41 68.29 ;
      RECT  50.17 71.88 51.32 72.02 ;
      RECT  49.76 70.97 50.33 71.3 ;
      RECT  50.97 68.95 52.59 69.12 ;
      RECT  50.59 69.18 50.76 69.36 ;
      RECT  52.3 68.89 52.59 68.95 ;
      RECT  50.53 68.89 50.82 69.18 ;
      RECT  50.81 71.38 51.1 71.44 ;
      RECT  50.81 71.15 51.1 71.21 ;
      RECT  52.04 68.59 52.33 68.67 ;
      RECT  52.29 70.44 52.58 70.5 ;
      RECT  50.17 71.86 51.04 71.88 ;
      RECT  51.76 70.44 52.11 70.53 ;
      RECT  52.29 74.71 52.58 74.65 ;
      RECT  52.04 76.54 52.33 76.48 ;
      RECT  49.61 76.48 52.69 76.33 ;
      RECT  50.06 72.75 50.41 72.4 ;
      RECT  50.81 73.71 52.0 73.54 ;
      RECT  52.3 75.8 52.59 75.74 ;
      RECT  50.17 73.62 50.33 73.06 ;
      RECT  51.76 74.74 52.11 74.65 ;
      RECT  50.97 75.8 51.32 75.71 ;
      RECT  50.97 76.06 51.32 75.97 ;
      RECT  50.59 75.56 51.04 75.42 ;
      RECT  51.77 73.04 52.06 72.75 ;
      RECT  51.76 74.65 52.58 74.48 ;
      RECT  51.03 72.9 51.32 72.75 ;
      RECT  51.83 73.54 52.0 73.04 ;
      RECT  50.87 75.42 51.04 73.77 ;
      RECT  50.06 76.98 50.41 76.63 ;
      RECT  50.17 73.04 51.32 72.9 ;
      RECT  49.76 73.95 50.33 73.62 ;
      RECT  50.97 75.97 52.59 75.8 ;
      RECT  50.59 75.74 50.76 75.56 ;
      RECT  52.3 76.03 52.59 75.97 ;
      RECT  50.53 76.03 50.82 75.74 ;
      RECT  50.81 73.54 51.1 73.48 ;
      RECT  50.81 73.77 51.1 73.71 ;
      RECT  52.04 76.33 52.33 76.25 ;
      RECT  52.29 74.48 52.58 74.42 ;
      RECT  50.17 73.06 51.04 73.04 ;
      RECT  51.76 74.48 52.11 74.39 ;
      RECT  52.29 78.91 52.58 78.97 ;
      RECT  52.04 77.08 52.33 77.14 ;
      RECT  49.61 77.14 52.69 77.29 ;
      RECT  50.06 80.87 50.41 81.22 ;
      RECT  50.81 79.91 52.0 80.08 ;
      RECT  52.3 77.82 52.59 77.88 ;
      RECT  50.17 80.0 50.33 80.56 ;
      RECT  51.76 78.88 52.11 78.97 ;
      RECT  50.97 77.82 51.32 77.91 ;
      RECT  50.97 77.56 51.32 77.65 ;
      RECT  50.59 78.06 51.04 78.2 ;
      RECT  51.77 80.58 52.06 80.87 ;
      RECT  51.76 78.97 52.58 79.14 ;
      RECT  51.03 80.72 51.32 80.87 ;
      RECT  51.83 80.08 52.0 80.58 ;
      RECT  50.87 78.2 51.04 79.85 ;
      RECT  50.06 76.64 50.41 76.99 ;
      RECT  50.17 80.58 51.32 80.72 ;
      RECT  49.76 79.67 50.33 80.0 ;
      RECT  50.97 77.65 52.59 77.82 ;
      RECT  50.59 77.88 50.76 78.06 ;
      RECT  52.3 77.59 52.59 77.65 ;
      RECT  50.53 77.59 50.82 77.88 ;
      RECT  50.81 80.08 51.1 80.14 ;
      RECT  50.81 79.85 51.1 79.91 ;
      RECT  52.04 77.29 52.33 77.37 ;
      RECT  52.29 79.14 52.58 79.2 ;
      RECT  50.17 80.56 51.04 80.58 ;
      RECT  51.76 79.14 52.11 79.23 ;
      RECT  52.29 83.41 52.58 83.35 ;
      RECT  52.04 85.24 52.33 85.18 ;
      RECT  49.61 85.18 52.69 85.03 ;
      RECT  50.06 81.45 50.41 81.1 ;
      RECT  50.81 82.41 52.0 82.24 ;
      RECT  52.3 84.5 52.59 84.44 ;
      RECT  50.17 82.32 50.33 81.76 ;
      RECT  51.76 83.44 52.11 83.35 ;
      RECT  50.97 84.5 51.32 84.41 ;
      RECT  50.97 84.76 51.32 84.67 ;
      RECT  50.59 84.26 51.04 84.12 ;
      RECT  51.77 81.74 52.06 81.45 ;
      RECT  51.76 83.35 52.58 83.18 ;
      RECT  51.03 81.6 51.32 81.45 ;
      RECT  51.83 82.24 52.0 81.74 ;
      RECT  50.87 84.12 51.04 82.47 ;
      RECT  50.06 85.68 50.41 85.33 ;
      RECT  50.17 81.74 51.32 81.6 ;
      RECT  49.76 82.65 50.33 82.32 ;
      RECT  50.97 84.67 52.59 84.5 ;
      RECT  50.59 84.44 50.76 84.26 ;
      RECT  52.3 84.73 52.59 84.67 ;
      RECT  50.53 84.73 50.82 84.44 ;
      RECT  50.81 82.24 51.1 82.18 ;
      RECT  50.81 82.47 51.1 82.41 ;
      RECT  52.04 85.03 52.33 84.95 ;
      RECT  52.29 83.18 52.58 83.12 ;
      RECT  50.17 81.76 51.04 81.74 ;
      RECT  51.76 83.18 52.11 83.09 ;
      RECT  52.29 87.61 52.58 87.67 ;
      RECT  52.04 85.78 52.33 85.84 ;
      RECT  49.61 85.84 52.69 85.99 ;
      RECT  50.06 89.57 50.41 89.92 ;
      RECT  50.81 88.61 52.0 88.78 ;
      RECT  52.3 86.52 52.59 86.58 ;
      RECT  50.17 88.7 50.33 89.26 ;
      RECT  51.76 87.58 52.11 87.67 ;
      RECT  50.97 86.52 51.32 86.61 ;
      RECT  50.97 86.26 51.32 86.35 ;
      RECT  50.59 86.76 51.04 86.9 ;
      RECT  51.77 89.28 52.06 89.57 ;
      RECT  51.76 87.67 52.58 87.84 ;
      RECT  51.03 89.42 51.32 89.57 ;
      RECT  51.83 88.78 52.0 89.28 ;
      RECT  50.87 86.9 51.04 88.55 ;
      RECT  50.06 85.34 50.41 85.69 ;
      RECT  50.17 89.28 51.32 89.42 ;
      RECT  49.76 88.37 50.33 88.7 ;
      RECT  50.97 86.35 52.59 86.52 ;
      RECT  50.59 86.58 50.76 86.76 ;
      RECT  52.3 86.29 52.59 86.35 ;
      RECT  50.53 86.29 50.82 86.58 ;
      RECT  50.81 88.78 51.1 88.84 ;
      RECT  50.81 88.55 51.1 88.61 ;
      RECT  52.04 85.99 52.33 86.07 ;
      RECT  52.29 87.84 52.58 87.9 ;
      RECT  50.17 89.26 51.04 89.28 ;
      RECT  51.76 87.84 52.11 87.93 ;
      RECT  52.29 92.11 52.58 92.05 ;
      RECT  52.04 93.94 52.33 93.88 ;
      RECT  49.61 93.88 52.69 93.73 ;
      RECT  50.06 90.15 50.41 89.8 ;
      RECT  50.81 91.11 52.0 90.94 ;
      RECT  52.3 93.2 52.59 93.14 ;
      RECT  50.17 91.02 50.33 90.46 ;
      RECT  51.76 92.14 52.11 92.05 ;
      RECT  50.97 93.2 51.32 93.11 ;
      RECT  50.97 93.46 51.32 93.37 ;
      RECT  50.59 92.96 51.04 92.82 ;
      RECT  51.77 90.44 52.06 90.15 ;
      RECT  51.76 92.05 52.58 91.88 ;
      RECT  51.03 90.3 51.32 90.15 ;
      RECT  51.83 90.94 52.0 90.44 ;
      RECT  50.87 92.82 51.04 91.17 ;
      RECT  50.06 94.38 50.41 94.03 ;
      RECT  50.17 90.44 51.32 90.3 ;
      RECT  49.76 91.35 50.33 91.02 ;
      RECT  50.97 93.37 52.59 93.2 ;
      RECT  50.59 93.14 50.76 92.96 ;
      RECT  52.3 93.43 52.59 93.37 ;
      RECT  50.53 93.43 50.82 93.14 ;
      RECT  50.81 90.94 51.1 90.88 ;
      RECT  50.81 91.17 51.1 91.11 ;
      RECT  52.04 93.73 52.33 93.65 ;
      RECT  52.29 91.88 52.58 91.82 ;
      RECT  50.17 90.46 51.04 90.44 ;
      RECT  51.76 91.88 52.11 91.79 ;
      RECT  52.29 96.31 52.58 96.37 ;
      RECT  52.04 94.48 52.33 94.54 ;
      RECT  49.61 94.54 52.69 94.69 ;
      RECT  50.06 98.27 50.41 98.62 ;
      RECT  50.81 97.31 52.0 97.48 ;
      RECT  52.3 95.22 52.59 95.28 ;
      RECT  50.17 97.4 50.33 97.96 ;
      RECT  51.76 96.28 52.11 96.37 ;
      RECT  50.97 95.22 51.32 95.31 ;
      RECT  50.97 94.96 51.32 95.05 ;
      RECT  50.59 95.46 51.04 95.6 ;
      RECT  51.77 97.98 52.06 98.27 ;
      RECT  51.76 96.37 52.58 96.54 ;
      RECT  51.03 98.12 51.32 98.27 ;
      RECT  51.83 97.48 52.0 97.98 ;
      RECT  50.87 95.6 51.04 97.25 ;
      RECT  50.06 94.04 50.41 94.39 ;
      RECT  50.17 97.98 51.32 98.12 ;
      RECT  49.76 97.07 50.33 97.4 ;
      RECT  50.97 95.05 52.59 95.22 ;
      RECT  50.59 95.28 50.76 95.46 ;
      RECT  52.3 94.99 52.59 95.05 ;
      RECT  50.53 94.99 50.82 95.28 ;
      RECT  50.81 97.48 51.1 97.54 ;
      RECT  50.81 97.25 51.1 97.31 ;
      RECT  52.04 94.69 52.33 94.77 ;
      RECT  52.29 96.54 52.58 96.6 ;
      RECT  50.17 97.96 51.04 97.98 ;
      RECT  51.76 96.54 52.11 96.63 ;
      RECT  52.29 100.81 52.58 100.75 ;
      RECT  52.04 102.64 52.33 102.58 ;
      RECT  49.61 102.58 52.69 102.43 ;
      RECT  50.06 98.85 50.41 98.5 ;
      RECT  50.81 99.81 52.0 99.64 ;
      RECT  52.3 101.9 52.59 101.84 ;
      RECT  50.17 99.72 50.33 99.16 ;
      RECT  51.76 100.84 52.11 100.75 ;
      RECT  50.97 101.9 51.32 101.81 ;
      RECT  50.97 102.16 51.32 102.07 ;
      RECT  50.59 101.66 51.04 101.52 ;
      RECT  51.77 99.14 52.06 98.85 ;
      RECT  51.76 100.75 52.58 100.58 ;
      RECT  51.03 99.0 51.32 98.85 ;
      RECT  51.83 99.64 52.0 99.14 ;
      RECT  50.87 101.52 51.04 99.87 ;
      RECT  50.06 103.08 50.41 102.73 ;
      RECT  50.17 99.14 51.32 99.0 ;
      RECT  49.76 100.05 50.33 99.72 ;
      RECT  50.97 102.07 52.59 101.9 ;
      RECT  50.59 101.84 50.76 101.66 ;
      RECT  52.3 102.13 52.59 102.07 ;
      RECT  50.53 102.13 50.82 101.84 ;
      RECT  50.81 99.64 51.1 99.58 ;
      RECT  50.81 99.87 51.1 99.81 ;
      RECT  52.04 102.43 52.33 102.35 ;
      RECT  52.29 100.58 52.58 100.52 ;
      RECT  50.17 99.16 51.04 99.14 ;
      RECT  51.76 100.58 52.11 100.49 ;
      RECT  55.37 35.41 55.66 35.47 ;
      RECT  55.12 33.58 55.41 33.64 ;
      RECT  52.69 33.64 55.77 33.79 ;
      RECT  53.14 37.37 53.49 37.72 ;
      RECT  53.89 36.41 55.08 36.58 ;
      RECT  55.38 34.32 55.67 34.38 ;
      RECT  53.25 36.5 53.41 37.06 ;
      RECT  54.84 35.38 55.19 35.47 ;
      RECT  54.05 34.32 54.4 34.41 ;
      RECT  54.05 34.06 54.4 34.15 ;
      RECT  53.67 34.56 54.12 34.7 ;
      RECT  54.85 37.08 55.14 37.37 ;
      RECT  54.84 35.47 55.66 35.64 ;
      RECT  54.11 37.22 54.4 37.37 ;
      RECT  54.91 36.58 55.08 37.08 ;
      RECT  53.95 34.7 54.12 36.35 ;
      RECT  53.14 33.14 53.49 33.49 ;
      RECT  53.25 37.08 54.4 37.22 ;
      RECT  52.84 36.17 53.41 36.5 ;
      RECT  54.05 34.15 55.67 34.32 ;
      RECT  53.67 34.38 53.84 34.56 ;
      RECT  55.38 34.09 55.67 34.15 ;
      RECT  53.61 34.09 53.9 34.38 ;
      RECT  53.89 36.58 54.18 36.64 ;
      RECT  53.89 36.35 54.18 36.41 ;
      RECT  55.12 33.79 55.41 33.87 ;
      RECT  55.37 35.64 55.66 35.7 ;
      RECT  53.25 37.06 54.12 37.08 ;
      RECT  54.84 35.64 55.19 35.73 ;
      RECT  55.37 39.91 55.66 39.85 ;
      RECT  55.12 41.74 55.41 41.68 ;
      RECT  52.69 41.68 55.77 41.53 ;
      RECT  53.14 37.95 53.49 37.6 ;
      RECT  53.89 38.91 55.08 38.74 ;
      RECT  55.38 41.0 55.67 40.94 ;
      RECT  53.25 38.82 53.41 38.26 ;
      RECT  54.84 39.94 55.19 39.85 ;
      RECT  54.05 41.0 54.4 40.91 ;
      RECT  54.05 41.26 54.4 41.17 ;
      RECT  53.67 40.76 54.12 40.62 ;
      RECT  54.85 38.24 55.14 37.95 ;
      RECT  54.84 39.85 55.66 39.68 ;
      RECT  54.11 38.1 54.4 37.95 ;
      RECT  54.91 38.74 55.08 38.24 ;
      RECT  53.95 40.62 54.12 38.97 ;
      RECT  53.14 42.18 53.49 41.83 ;
      RECT  53.25 38.24 54.4 38.1 ;
      RECT  52.84 39.15 53.41 38.82 ;
      RECT  54.05 41.17 55.67 41.0 ;
      RECT  53.67 40.94 53.84 40.76 ;
      RECT  55.38 41.23 55.67 41.17 ;
      RECT  53.61 41.23 53.9 40.94 ;
      RECT  53.89 38.74 54.18 38.68 ;
      RECT  53.89 38.97 54.18 38.91 ;
      RECT  55.12 41.53 55.41 41.45 ;
      RECT  55.37 39.68 55.66 39.62 ;
      RECT  53.25 38.26 54.12 38.24 ;
      RECT  54.84 39.68 55.19 39.59 ;
      RECT  55.37 44.11 55.66 44.17 ;
      RECT  55.12 42.28 55.41 42.34 ;
      RECT  52.69 42.34 55.77 42.49 ;
      RECT  53.14 46.07 53.49 46.42 ;
      RECT  53.89 45.11 55.08 45.28 ;
      RECT  55.38 43.02 55.67 43.08 ;
      RECT  53.25 45.2 53.41 45.76 ;
      RECT  54.84 44.08 55.19 44.17 ;
      RECT  54.05 43.02 54.4 43.11 ;
      RECT  54.05 42.76 54.4 42.85 ;
      RECT  53.67 43.26 54.12 43.4 ;
      RECT  54.85 45.78 55.14 46.07 ;
      RECT  54.84 44.17 55.66 44.34 ;
      RECT  54.11 45.92 54.4 46.07 ;
      RECT  54.91 45.28 55.08 45.78 ;
      RECT  53.95 43.4 54.12 45.05 ;
      RECT  53.14 41.84 53.49 42.19 ;
      RECT  53.25 45.78 54.4 45.92 ;
      RECT  52.84 44.87 53.41 45.2 ;
      RECT  54.05 42.85 55.67 43.02 ;
      RECT  53.67 43.08 53.84 43.26 ;
      RECT  55.38 42.79 55.67 42.85 ;
      RECT  53.61 42.79 53.9 43.08 ;
      RECT  53.89 45.28 54.18 45.34 ;
      RECT  53.89 45.05 54.18 45.11 ;
      RECT  55.12 42.49 55.41 42.57 ;
      RECT  55.37 44.34 55.66 44.4 ;
      RECT  53.25 45.76 54.12 45.78 ;
      RECT  54.84 44.34 55.19 44.43 ;
      RECT  55.37 48.61 55.66 48.55 ;
      RECT  55.12 50.44 55.41 50.38 ;
      RECT  52.69 50.38 55.77 50.23 ;
      RECT  53.14 46.65 53.49 46.3 ;
      RECT  53.89 47.61 55.08 47.44 ;
      RECT  55.38 49.7 55.67 49.64 ;
      RECT  53.25 47.52 53.41 46.96 ;
      RECT  54.84 48.64 55.19 48.55 ;
      RECT  54.05 49.7 54.4 49.61 ;
      RECT  54.05 49.96 54.4 49.87 ;
      RECT  53.67 49.46 54.12 49.32 ;
      RECT  54.85 46.94 55.14 46.65 ;
      RECT  54.84 48.55 55.66 48.38 ;
      RECT  54.11 46.8 54.4 46.65 ;
      RECT  54.91 47.44 55.08 46.94 ;
      RECT  53.95 49.32 54.12 47.67 ;
      RECT  53.14 50.88 53.49 50.53 ;
      RECT  53.25 46.94 54.4 46.8 ;
      RECT  52.84 47.85 53.41 47.52 ;
      RECT  54.05 49.87 55.67 49.7 ;
      RECT  53.67 49.64 53.84 49.46 ;
      RECT  55.38 49.93 55.67 49.87 ;
      RECT  53.61 49.93 53.9 49.64 ;
      RECT  53.89 47.44 54.18 47.38 ;
      RECT  53.89 47.67 54.18 47.61 ;
      RECT  55.12 50.23 55.41 50.15 ;
      RECT  55.37 48.38 55.66 48.32 ;
      RECT  53.25 46.96 54.12 46.94 ;
      RECT  54.84 48.38 55.19 48.29 ;
      RECT  55.37 52.81 55.66 52.87 ;
      RECT  55.12 50.98 55.41 51.04 ;
      RECT  52.69 51.04 55.77 51.19 ;
      RECT  53.14 54.77 53.49 55.12 ;
      RECT  53.89 53.81 55.08 53.98 ;
      RECT  55.38 51.72 55.67 51.78 ;
      RECT  53.25 53.9 53.41 54.46 ;
      RECT  54.84 52.78 55.19 52.87 ;
      RECT  54.05 51.72 54.4 51.81 ;
      RECT  54.05 51.46 54.4 51.55 ;
      RECT  53.67 51.96 54.12 52.1 ;
      RECT  54.85 54.48 55.14 54.77 ;
      RECT  54.84 52.87 55.66 53.04 ;
      RECT  54.11 54.62 54.4 54.77 ;
      RECT  54.91 53.98 55.08 54.48 ;
      RECT  53.95 52.1 54.12 53.75 ;
      RECT  53.14 50.54 53.49 50.89 ;
      RECT  53.25 54.48 54.4 54.62 ;
      RECT  52.84 53.57 53.41 53.9 ;
      RECT  54.05 51.55 55.67 51.72 ;
      RECT  53.67 51.78 53.84 51.96 ;
      RECT  55.38 51.49 55.67 51.55 ;
      RECT  53.61 51.49 53.9 51.78 ;
      RECT  53.89 53.98 54.18 54.04 ;
      RECT  53.89 53.75 54.18 53.81 ;
      RECT  55.12 51.19 55.41 51.27 ;
      RECT  55.37 53.04 55.66 53.1 ;
      RECT  53.25 54.46 54.12 54.48 ;
      RECT  54.84 53.04 55.19 53.13 ;
      RECT  55.37 57.31 55.66 57.25 ;
      RECT  55.12 59.14 55.41 59.08 ;
      RECT  52.69 59.08 55.77 58.93 ;
      RECT  53.14 55.35 53.49 55.0 ;
      RECT  53.89 56.31 55.08 56.14 ;
      RECT  55.38 58.4 55.67 58.34 ;
      RECT  53.25 56.22 53.41 55.66 ;
      RECT  54.84 57.34 55.19 57.25 ;
      RECT  54.05 58.4 54.4 58.31 ;
      RECT  54.05 58.66 54.4 58.57 ;
      RECT  53.67 58.16 54.12 58.02 ;
      RECT  54.85 55.64 55.14 55.35 ;
      RECT  54.84 57.25 55.66 57.08 ;
      RECT  54.11 55.5 54.4 55.35 ;
      RECT  54.91 56.14 55.08 55.64 ;
      RECT  53.95 58.02 54.12 56.37 ;
      RECT  53.14 59.58 53.49 59.23 ;
      RECT  53.25 55.64 54.4 55.5 ;
      RECT  52.84 56.55 53.41 56.22 ;
      RECT  54.05 58.57 55.67 58.4 ;
      RECT  53.67 58.34 53.84 58.16 ;
      RECT  55.38 58.63 55.67 58.57 ;
      RECT  53.61 58.63 53.9 58.34 ;
      RECT  53.89 56.14 54.18 56.08 ;
      RECT  53.89 56.37 54.18 56.31 ;
      RECT  55.12 58.93 55.41 58.85 ;
      RECT  55.37 57.08 55.66 57.02 ;
      RECT  53.25 55.66 54.12 55.64 ;
      RECT  54.84 57.08 55.19 56.99 ;
      RECT  55.37 61.51 55.66 61.57 ;
      RECT  55.12 59.68 55.41 59.74 ;
      RECT  52.69 59.74 55.77 59.89 ;
      RECT  53.14 63.47 53.49 63.82 ;
      RECT  53.89 62.51 55.08 62.68 ;
      RECT  55.38 60.42 55.67 60.48 ;
      RECT  53.25 62.6 53.41 63.16 ;
      RECT  54.84 61.48 55.19 61.57 ;
      RECT  54.05 60.42 54.4 60.51 ;
      RECT  54.05 60.16 54.4 60.25 ;
      RECT  53.67 60.66 54.12 60.8 ;
      RECT  54.85 63.18 55.14 63.47 ;
      RECT  54.84 61.57 55.66 61.74 ;
      RECT  54.11 63.32 54.4 63.47 ;
      RECT  54.91 62.68 55.08 63.18 ;
      RECT  53.95 60.8 54.12 62.45 ;
      RECT  53.14 59.24 53.49 59.59 ;
      RECT  53.25 63.18 54.4 63.32 ;
      RECT  52.84 62.27 53.41 62.6 ;
      RECT  54.05 60.25 55.67 60.42 ;
      RECT  53.67 60.48 53.84 60.66 ;
      RECT  55.38 60.19 55.67 60.25 ;
      RECT  53.61 60.19 53.9 60.48 ;
      RECT  53.89 62.68 54.18 62.74 ;
      RECT  53.89 62.45 54.18 62.51 ;
      RECT  55.12 59.89 55.41 59.97 ;
      RECT  55.37 61.74 55.66 61.8 ;
      RECT  53.25 63.16 54.12 63.18 ;
      RECT  54.84 61.74 55.19 61.83 ;
      RECT  55.37 66.01 55.66 65.95 ;
      RECT  55.12 67.84 55.41 67.78 ;
      RECT  52.69 67.78 55.77 67.63 ;
      RECT  53.14 64.05 53.49 63.7 ;
      RECT  53.89 65.01 55.08 64.84 ;
      RECT  55.38 67.1 55.67 67.04 ;
      RECT  53.25 64.92 53.41 64.36 ;
      RECT  54.84 66.04 55.19 65.95 ;
      RECT  54.05 67.1 54.4 67.01 ;
      RECT  54.05 67.36 54.4 67.27 ;
      RECT  53.67 66.86 54.12 66.72 ;
      RECT  54.85 64.34 55.14 64.05 ;
      RECT  54.84 65.95 55.66 65.78 ;
      RECT  54.11 64.2 54.4 64.05 ;
      RECT  54.91 64.84 55.08 64.34 ;
      RECT  53.95 66.72 54.12 65.07 ;
      RECT  53.14 68.28 53.49 67.93 ;
      RECT  53.25 64.34 54.4 64.2 ;
      RECT  52.84 65.25 53.41 64.92 ;
      RECT  54.05 67.27 55.67 67.1 ;
      RECT  53.67 67.04 53.84 66.86 ;
      RECT  55.38 67.33 55.67 67.27 ;
      RECT  53.61 67.33 53.9 67.04 ;
      RECT  53.89 64.84 54.18 64.78 ;
      RECT  53.89 65.07 54.18 65.01 ;
      RECT  55.12 67.63 55.41 67.55 ;
      RECT  55.37 65.78 55.66 65.72 ;
      RECT  53.25 64.36 54.12 64.34 ;
      RECT  54.84 65.78 55.19 65.69 ;
      RECT  55.37 70.21 55.66 70.27 ;
      RECT  55.12 68.38 55.41 68.44 ;
      RECT  52.69 68.44 55.77 68.59 ;
      RECT  53.14 72.17 53.49 72.52 ;
      RECT  53.89 71.21 55.08 71.38 ;
      RECT  55.38 69.12 55.67 69.18 ;
      RECT  53.25 71.3 53.41 71.86 ;
      RECT  54.84 70.18 55.19 70.27 ;
      RECT  54.05 69.12 54.4 69.21 ;
      RECT  54.05 68.86 54.4 68.95 ;
      RECT  53.67 69.36 54.12 69.5 ;
      RECT  54.85 71.88 55.14 72.17 ;
      RECT  54.84 70.27 55.66 70.44 ;
      RECT  54.11 72.02 54.4 72.17 ;
      RECT  54.91 71.38 55.08 71.88 ;
      RECT  53.95 69.5 54.12 71.15 ;
      RECT  53.14 67.94 53.49 68.29 ;
      RECT  53.25 71.88 54.4 72.02 ;
      RECT  52.84 70.97 53.41 71.3 ;
      RECT  54.05 68.95 55.67 69.12 ;
      RECT  53.67 69.18 53.84 69.36 ;
      RECT  55.38 68.89 55.67 68.95 ;
      RECT  53.61 68.89 53.9 69.18 ;
      RECT  53.89 71.38 54.18 71.44 ;
      RECT  53.89 71.15 54.18 71.21 ;
      RECT  55.12 68.59 55.41 68.67 ;
      RECT  55.37 70.44 55.66 70.5 ;
      RECT  53.25 71.86 54.12 71.88 ;
      RECT  54.84 70.44 55.19 70.53 ;
      RECT  55.37 74.71 55.66 74.65 ;
      RECT  55.12 76.54 55.41 76.48 ;
      RECT  52.69 76.48 55.77 76.33 ;
      RECT  53.14 72.75 53.49 72.4 ;
      RECT  53.89 73.71 55.08 73.54 ;
      RECT  55.38 75.8 55.67 75.74 ;
      RECT  53.25 73.62 53.41 73.06 ;
      RECT  54.84 74.74 55.19 74.65 ;
      RECT  54.05 75.8 54.4 75.71 ;
      RECT  54.05 76.06 54.4 75.97 ;
      RECT  53.67 75.56 54.12 75.42 ;
      RECT  54.85 73.04 55.14 72.75 ;
      RECT  54.84 74.65 55.66 74.48 ;
      RECT  54.11 72.9 54.4 72.75 ;
      RECT  54.91 73.54 55.08 73.04 ;
      RECT  53.95 75.42 54.12 73.77 ;
      RECT  53.14 76.98 53.49 76.63 ;
      RECT  53.25 73.04 54.4 72.9 ;
      RECT  52.84 73.95 53.41 73.62 ;
      RECT  54.05 75.97 55.67 75.8 ;
      RECT  53.67 75.74 53.84 75.56 ;
      RECT  55.38 76.03 55.67 75.97 ;
      RECT  53.61 76.03 53.9 75.74 ;
      RECT  53.89 73.54 54.18 73.48 ;
      RECT  53.89 73.77 54.18 73.71 ;
      RECT  55.12 76.33 55.41 76.25 ;
      RECT  55.37 74.48 55.66 74.42 ;
      RECT  53.25 73.06 54.12 73.04 ;
      RECT  54.84 74.48 55.19 74.39 ;
      RECT  55.37 78.91 55.66 78.97 ;
      RECT  55.12 77.08 55.41 77.14 ;
      RECT  52.69 77.14 55.77 77.29 ;
      RECT  53.14 80.87 53.49 81.22 ;
      RECT  53.89 79.91 55.08 80.08 ;
      RECT  55.38 77.82 55.67 77.88 ;
      RECT  53.25 80.0 53.41 80.56 ;
      RECT  54.84 78.88 55.19 78.97 ;
      RECT  54.05 77.82 54.4 77.91 ;
      RECT  54.05 77.56 54.4 77.65 ;
      RECT  53.67 78.06 54.12 78.2 ;
      RECT  54.85 80.58 55.14 80.87 ;
      RECT  54.84 78.97 55.66 79.14 ;
      RECT  54.11 80.72 54.4 80.87 ;
      RECT  54.91 80.08 55.08 80.58 ;
      RECT  53.95 78.2 54.12 79.85 ;
      RECT  53.14 76.64 53.49 76.99 ;
      RECT  53.25 80.58 54.4 80.72 ;
      RECT  52.84 79.67 53.41 80.0 ;
      RECT  54.05 77.65 55.67 77.82 ;
      RECT  53.67 77.88 53.84 78.06 ;
      RECT  55.38 77.59 55.67 77.65 ;
      RECT  53.61 77.59 53.9 77.88 ;
      RECT  53.89 80.08 54.18 80.14 ;
      RECT  53.89 79.85 54.18 79.91 ;
      RECT  55.12 77.29 55.41 77.37 ;
      RECT  55.37 79.14 55.66 79.2 ;
      RECT  53.25 80.56 54.12 80.58 ;
      RECT  54.84 79.14 55.19 79.23 ;
      RECT  55.37 83.41 55.66 83.35 ;
      RECT  55.12 85.24 55.41 85.18 ;
      RECT  52.69 85.18 55.77 85.03 ;
      RECT  53.14 81.45 53.49 81.1 ;
      RECT  53.89 82.41 55.08 82.24 ;
      RECT  55.38 84.5 55.67 84.44 ;
      RECT  53.25 82.32 53.41 81.76 ;
      RECT  54.84 83.44 55.19 83.35 ;
      RECT  54.05 84.5 54.4 84.41 ;
      RECT  54.05 84.76 54.4 84.67 ;
      RECT  53.67 84.26 54.12 84.12 ;
      RECT  54.85 81.74 55.14 81.45 ;
      RECT  54.84 83.35 55.66 83.18 ;
      RECT  54.11 81.6 54.4 81.45 ;
      RECT  54.91 82.24 55.08 81.74 ;
      RECT  53.95 84.12 54.12 82.47 ;
      RECT  53.14 85.68 53.49 85.33 ;
      RECT  53.25 81.74 54.4 81.6 ;
      RECT  52.84 82.65 53.41 82.32 ;
      RECT  54.05 84.67 55.67 84.5 ;
      RECT  53.67 84.44 53.84 84.26 ;
      RECT  55.38 84.73 55.67 84.67 ;
      RECT  53.61 84.73 53.9 84.44 ;
      RECT  53.89 82.24 54.18 82.18 ;
      RECT  53.89 82.47 54.18 82.41 ;
      RECT  55.12 85.03 55.41 84.95 ;
      RECT  55.37 83.18 55.66 83.12 ;
      RECT  53.25 81.76 54.12 81.74 ;
      RECT  54.84 83.18 55.19 83.09 ;
      RECT  55.37 87.61 55.66 87.67 ;
      RECT  55.12 85.78 55.41 85.84 ;
      RECT  52.69 85.84 55.77 85.99 ;
      RECT  53.14 89.57 53.49 89.92 ;
      RECT  53.89 88.61 55.08 88.78 ;
      RECT  55.38 86.52 55.67 86.58 ;
      RECT  53.25 88.7 53.41 89.26 ;
      RECT  54.84 87.58 55.19 87.67 ;
      RECT  54.05 86.52 54.4 86.61 ;
      RECT  54.05 86.26 54.4 86.35 ;
      RECT  53.67 86.76 54.12 86.9 ;
      RECT  54.85 89.28 55.14 89.57 ;
      RECT  54.84 87.67 55.66 87.84 ;
      RECT  54.11 89.42 54.4 89.57 ;
      RECT  54.91 88.78 55.08 89.28 ;
      RECT  53.95 86.9 54.12 88.55 ;
      RECT  53.14 85.34 53.49 85.69 ;
      RECT  53.25 89.28 54.4 89.42 ;
      RECT  52.84 88.37 53.41 88.7 ;
      RECT  54.05 86.35 55.67 86.52 ;
      RECT  53.67 86.58 53.84 86.76 ;
      RECT  55.38 86.29 55.67 86.35 ;
      RECT  53.61 86.29 53.9 86.58 ;
      RECT  53.89 88.78 54.18 88.84 ;
      RECT  53.89 88.55 54.18 88.61 ;
      RECT  55.12 85.99 55.41 86.07 ;
      RECT  55.37 87.84 55.66 87.9 ;
      RECT  53.25 89.26 54.12 89.28 ;
      RECT  54.84 87.84 55.19 87.93 ;
      RECT  55.37 92.11 55.66 92.05 ;
      RECT  55.12 93.94 55.41 93.88 ;
      RECT  52.69 93.88 55.77 93.73 ;
      RECT  53.14 90.15 53.49 89.8 ;
      RECT  53.89 91.11 55.08 90.94 ;
      RECT  55.38 93.2 55.67 93.14 ;
      RECT  53.25 91.02 53.41 90.46 ;
      RECT  54.84 92.14 55.19 92.05 ;
      RECT  54.05 93.2 54.4 93.11 ;
      RECT  54.05 93.46 54.4 93.37 ;
      RECT  53.67 92.96 54.12 92.82 ;
      RECT  54.85 90.44 55.14 90.15 ;
      RECT  54.84 92.05 55.66 91.88 ;
      RECT  54.11 90.3 54.4 90.15 ;
      RECT  54.91 90.94 55.08 90.44 ;
      RECT  53.95 92.82 54.12 91.17 ;
      RECT  53.14 94.38 53.49 94.03 ;
      RECT  53.25 90.44 54.4 90.3 ;
      RECT  52.84 91.35 53.41 91.02 ;
      RECT  54.05 93.37 55.67 93.2 ;
      RECT  53.67 93.14 53.84 92.96 ;
      RECT  55.38 93.43 55.67 93.37 ;
      RECT  53.61 93.43 53.9 93.14 ;
      RECT  53.89 90.94 54.18 90.88 ;
      RECT  53.89 91.17 54.18 91.11 ;
      RECT  55.12 93.73 55.41 93.65 ;
      RECT  55.37 91.88 55.66 91.82 ;
      RECT  53.25 90.46 54.12 90.44 ;
      RECT  54.84 91.88 55.19 91.79 ;
      RECT  55.37 96.31 55.66 96.37 ;
      RECT  55.12 94.48 55.41 94.54 ;
      RECT  52.69 94.54 55.77 94.69 ;
      RECT  53.14 98.27 53.49 98.62 ;
      RECT  53.89 97.31 55.08 97.48 ;
      RECT  55.38 95.22 55.67 95.28 ;
      RECT  53.25 97.4 53.41 97.96 ;
      RECT  54.84 96.28 55.19 96.37 ;
      RECT  54.05 95.22 54.4 95.31 ;
      RECT  54.05 94.96 54.4 95.05 ;
      RECT  53.67 95.46 54.12 95.6 ;
      RECT  54.85 97.98 55.14 98.27 ;
      RECT  54.84 96.37 55.66 96.54 ;
      RECT  54.11 98.12 54.4 98.27 ;
      RECT  54.91 97.48 55.08 97.98 ;
      RECT  53.95 95.6 54.12 97.25 ;
      RECT  53.14 94.04 53.49 94.39 ;
      RECT  53.25 97.98 54.4 98.12 ;
      RECT  52.84 97.07 53.41 97.4 ;
      RECT  54.05 95.05 55.67 95.22 ;
      RECT  53.67 95.28 53.84 95.46 ;
      RECT  55.38 94.99 55.67 95.05 ;
      RECT  53.61 94.99 53.9 95.28 ;
      RECT  53.89 97.48 54.18 97.54 ;
      RECT  53.89 97.25 54.18 97.31 ;
      RECT  55.12 94.69 55.41 94.77 ;
      RECT  55.37 96.54 55.66 96.6 ;
      RECT  53.25 97.96 54.12 97.98 ;
      RECT  54.84 96.54 55.19 96.63 ;
      RECT  55.37 100.81 55.66 100.75 ;
      RECT  55.12 102.64 55.41 102.58 ;
      RECT  52.69 102.58 55.77 102.43 ;
      RECT  53.14 98.85 53.49 98.5 ;
      RECT  53.89 99.81 55.08 99.64 ;
      RECT  55.38 101.9 55.67 101.84 ;
      RECT  53.25 99.72 53.41 99.16 ;
      RECT  54.84 100.84 55.19 100.75 ;
      RECT  54.05 101.9 54.4 101.81 ;
      RECT  54.05 102.16 54.4 102.07 ;
      RECT  53.67 101.66 54.12 101.52 ;
      RECT  54.85 99.14 55.14 98.85 ;
      RECT  54.84 100.75 55.66 100.58 ;
      RECT  54.11 99.0 54.4 98.85 ;
      RECT  54.91 99.64 55.08 99.14 ;
      RECT  53.95 101.52 54.12 99.87 ;
      RECT  53.14 103.08 53.49 102.73 ;
      RECT  53.25 99.14 54.4 99.0 ;
      RECT  52.84 100.05 53.41 99.72 ;
      RECT  54.05 102.07 55.67 101.9 ;
      RECT  53.67 101.84 53.84 101.66 ;
      RECT  55.38 102.13 55.67 102.07 ;
      RECT  53.61 102.13 53.9 101.84 ;
      RECT  53.89 99.64 54.18 99.58 ;
      RECT  53.89 99.87 54.18 99.81 ;
      RECT  55.12 102.43 55.41 102.35 ;
      RECT  55.37 100.58 55.66 100.52 ;
      RECT  53.25 99.16 54.12 99.14 ;
      RECT  54.84 100.58 55.19 100.49 ;
      RECT  49.61 33.64 55.77 33.79 ;
      RECT  49.61 41.53 55.77 41.68 ;
      RECT  49.61 42.34 55.77 42.49 ;
      RECT  49.61 50.23 55.77 50.38 ;
      RECT  49.61 51.04 55.77 51.19 ;
      RECT  49.61 58.93 55.77 59.08 ;
      RECT  49.61 59.74 55.77 59.89 ;
      RECT  49.61 67.63 55.77 67.78 ;
      RECT  49.61 68.44 55.77 68.59 ;
      RECT  49.61 76.33 55.77 76.48 ;
      RECT  49.61 77.14 55.77 77.29 ;
      RECT  49.61 85.03 55.77 85.18 ;
      RECT  49.61 85.84 55.77 85.99 ;
      RECT  49.61 93.73 55.77 93.88 ;
      RECT  49.61 94.54 55.77 94.69 ;
      RECT  49.61 102.43 55.77 102.58 ;
      RECT  49.21 26.71 49.5 26.77 ;
      RECT  48.96 24.88 49.25 24.94 ;
      RECT  46.53 24.94 49.61 25.09 ;
      RECT  46.98 28.67 47.33 29.02 ;
      RECT  47.73 27.71 48.92 27.88 ;
      RECT  49.22 25.62 49.51 25.68 ;
      RECT  47.09 27.8 47.25 28.36 ;
      RECT  48.68 26.68 49.03 26.77 ;
      RECT  47.89 25.62 48.24 25.71 ;
      RECT  47.89 25.36 48.24 25.45 ;
      RECT  47.51 25.86 47.96 26.0 ;
      RECT  48.69 28.38 48.98 28.67 ;
      RECT  48.68 26.77 49.5 26.94 ;
      RECT  47.95 28.52 48.24 28.67 ;
      RECT  48.75 27.88 48.92 28.38 ;
      RECT  47.79 26.0 47.96 27.65 ;
      RECT  46.98 24.44 47.33 24.79 ;
      RECT  47.09 28.38 48.24 28.52 ;
      RECT  46.68 27.47 47.25 27.8 ;
      RECT  47.89 25.45 49.51 25.62 ;
      RECT  47.51 25.68 47.68 25.86 ;
      RECT  49.22 25.39 49.51 25.45 ;
      RECT  47.45 25.39 47.74 25.68 ;
      RECT  47.73 27.88 48.02 27.94 ;
      RECT  47.73 27.65 48.02 27.71 ;
      RECT  48.96 25.09 49.25 25.17 ;
      RECT  49.21 26.94 49.5 27.0 ;
      RECT  47.09 28.36 47.96 28.38 ;
      RECT  48.68 26.94 49.03 27.03 ;
      RECT  49.21 31.21 49.5 31.15 ;
      RECT  48.96 33.04 49.25 32.98 ;
      RECT  46.53 32.98 49.61 32.83 ;
      RECT  46.98 29.25 47.33 28.9 ;
      RECT  47.73 30.21 48.92 30.04 ;
      RECT  49.22 32.3 49.51 32.24 ;
      RECT  47.09 30.12 47.25 29.56 ;
      RECT  48.68 31.24 49.03 31.15 ;
      RECT  47.89 32.3 48.24 32.21 ;
      RECT  47.89 32.56 48.24 32.47 ;
      RECT  47.51 32.06 47.96 31.92 ;
      RECT  48.69 29.54 48.98 29.25 ;
      RECT  48.68 31.15 49.5 30.98 ;
      RECT  47.95 29.4 48.24 29.25 ;
      RECT  48.75 30.04 48.92 29.54 ;
      RECT  47.79 31.92 47.96 30.27 ;
      RECT  46.98 33.48 47.33 33.13 ;
      RECT  47.09 29.54 48.24 29.4 ;
      RECT  46.68 30.45 47.25 30.12 ;
      RECT  47.89 32.47 49.51 32.3 ;
      RECT  47.51 32.24 47.68 32.06 ;
      RECT  49.22 32.53 49.51 32.47 ;
      RECT  47.45 32.53 47.74 32.24 ;
      RECT  47.73 30.04 48.02 29.98 ;
      RECT  47.73 30.27 48.02 30.21 ;
      RECT  48.96 32.83 49.25 32.75 ;
      RECT  49.21 30.98 49.5 30.92 ;
      RECT  47.09 29.56 47.96 29.54 ;
      RECT  48.68 30.98 49.03 30.89 ;
      RECT  49.21 35.41 49.5 35.47 ;
      RECT  48.96 33.58 49.25 33.64 ;
      RECT  46.53 33.64 49.61 33.79 ;
      RECT  46.98 37.37 47.33 37.72 ;
      RECT  47.73 36.41 48.92 36.58 ;
      RECT  49.22 34.32 49.51 34.38 ;
      RECT  47.09 36.5 47.25 37.06 ;
      RECT  48.68 35.38 49.03 35.47 ;
      RECT  47.89 34.32 48.24 34.41 ;
      RECT  47.89 34.06 48.24 34.15 ;
      RECT  47.51 34.56 47.96 34.7 ;
      RECT  48.69 37.08 48.98 37.37 ;
      RECT  48.68 35.47 49.5 35.64 ;
      RECT  47.95 37.22 48.24 37.37 ;
      RECT  48.75 36.58 48.92 37.08 ;
      RECT  47.79 34.7 47.96 36.35 ;
      RECT  46.98 33.14 47.33 33.49 ;
      RECT  47.09 37.08 48.24 37.22 ;
      RECT  46.68 36.17 47.25 36.5 ;
      RECT  47.89 34.15 49.51 34.32 ;
      RECT  47.51 34.38 47.68 34.56 ;
      RECT  49.22 34.09 49.51 34.15 ;
      RECT  47.45 34.09 47.74 34.38 ;
      RECT  47.73 36.58 48.02 36.64 ;
      RECT  47.73 36.35 48.02 36.41 ;
      RECT  48.96 33.79 49.25 33.87 ;
      RECT  49.21 35.64 49.5 35.7 ;
      RECT  47.09 37.06 47.96 37.08 ;
      RECT  48.68 35.64 49.03 35.73 ;
      RECT  49.21 39.91 49.5 39.85 ;
      RECT  48.96 41.74 49.25 41.68 ;
      RECT  46.53 41.68 49.61 41.53 ;
      RECT  46.98 37.95 47.33 37.6 ;
      RECT  47.73 38.91 48.92 38.74 ;
      RECT  49.22 41.0 49.51 40.94 ;
      RECT  47.09 38.82 47.25 38.26 ;
      RECT  48.68 39.94 49.03 39.85 ;
      RECT  47.89 41.0 48.24 40.91 ;
      RECT  47.89 41.26 48.24 41.17 ;
      RECT  47.51 40.76 47.96 40.62 ;
      RECT  48.69 38.24 48.98 37.95 ;
      RECT  48.68 39.85 49.5 39.68 ;
      RECT  47.95 38.1 48.24 37.95 ;
      RECT  48.75 38.74 48.92 38.24 ;
      RECT  47.79 40.62 47.96 38.97 ;
      RECT  46.98 42.18 47.33 41.83 ;
      RECT  47.09 38.24 48.24 38.1 ;
      RECT  46.68 39.15 47.25 38.82 ;
      RECT  47.89 41.17 49.51 41.0 ;
      RECT  47.51 40.94 47.68 40.76 ;
      RECT  49.22 41.23 49.51 41.17 ;
      RECT  47.45 41.23 47.74 40.94 ;
      RECT  47.73 38.74 48.02 38.68 ;
      RECT  47.73 38.97 48.02 38.91 ;
      RECT  48.96 41.53 49.25 41.45 ;
      RECT  49.21 39.68 49.5 39.62 ;
      RECT  47.09 38.26 47.96 38.24 ;
      RECT  48.68 39.68 49.03 39.59 ;
      RECT  49.21 44.11 49.5 44.17 ;
      RECT  48.96 42.28 49.25 42.34 ;
      RECT  46.53 42.34 49.61 42.49 ;
      RECT  46.98 46.07 47.33 46.42 ;
      RECT  47.73 45.11 48.92 45.28 ;
      RECT  49.22 43.02 49.51 43.08 ;
      RECT  47.09 45.2 47.25 45.76 ;
      RECT  48.68 44.08 49.03 44.17 ;
      RECT  47.89 43.02 48.24 43.11 ;
      RECT  47.89 42.76 48.24 42.85 ;
      RECT  47.51 43.26 47.96 43.4 ;
      RECT  48.69 45.78 48.98 46.07 ;
      RECT  48.68 44.17 49.5 44.34 ;
      RECT  47.95 45.92 48.24 46.07 ;
      RECT  48.75 45.28 48.92 45.78 ;
      RECT  47.79 43.4 47.96 45.05 ;
      RECT  46.98 41.84 47.33 42.19 ;
      RECT  47.09 45.78 48.24 45.92 ;
      RECT  46.68 44.87 47.25 45.2 ;
      RECT  47.89 42.85 49.51 43.02 ;
      RECT  47.51 43.08 47.68 43.26 ;
      RECT  49.22 42.79 49.51 42.85 ;
      RECT  47.45 42.79 47.74 43.08 ;
      RECT  47.73 45.28 48.02 45.34 ;
      RECT  47.73 45.05 48.02 45.11 ;
      RECT  48.96 42.49 49.25 42.57 ;
      RECT  49.21 44.34 49.5 44.4 ;
      RECT  47.09 45.76 47.96 45.78 ;
      RECT  48.68 44.34 49.03 44.43 ;
      RECT  49.21 48.61 49.5 48.55 ;
      RECT  48.96 50.44 49.25 50.38 ;
      RECT  46.53 50.38 49.61 50.23 ;
      RECT  46.98 46.65 47.33 46.3 ;
      RECT  47.73 47.61 48.92 47.44 ;
      RECT  49.22 49.7 49.51 49.64 ;
      RECT  47.09 47.52 47.25 46.96 ;
      RECT  48.68 48.64 49.03 48.55 ;
      RECT  47.89 49.7 48.24 49.61 ;
      RECT  47.89 49.96 48.24 49.87 ;
      RECT  47.51 49.46 47.96 49.32 ;
      RECT  48.69 46.94 48.98 46.65 ;
      RECT  48.68 48.55 49.5 48.38 ;
      RECT  47.95 46.8 48.24 46.65 ;
      RECT  48.75 47.44 48.92 46.94 ;
      RECT  47.79 49.32 47.96 47.67 ;
      RECT  46.98 50.88 47.33 50.53 ;
      RECT  47.09 46.94 48.24 46.8 ;
      RECT  46.68 47.85 47.25 47.52 ;
      RECT  47.89 49.87 49.51 49.7 ;
      RECT  47.51 49.64 47.68 49.46 ;
      RECT  49.22 49.93 49.51 49.87 ;
      RECT  47.45 49.93 47.74 49.64 ;
      RECT  47.73 47.44 48.02 47.38 ;
      RECT  47.73 47.67 48.02 47.61 ;
      RECT  48.96 50.23 49.25 50.15 ;
      RECT  49.21 48.38 49.5 48.32 ;
      RECT  47.09 46.96 47.96 46.94 ;
      RECT  48.68 48.38 49.03 48.29 ;
      RECT  49.21 52.81 49.5 52.87 ;
      RECT  48.96 50.98 49.25 51.04 ;
      RECT  46.53 51.04 49.61 51.19 ;
      RECT  46.98 54.77 47.33 55.12 ;
      RECT  47.73 53.81 48.92 53.98 ;
      RECT  49.22 51.72 49.51 51.78 ;
      RECT  47.09 53.9 47.25 54.46 ;
      RECT  48.68 52.78 49.03 52.87 ;
      RECT  47.89 51.72 48.24 51.81 ;
      RECT  47.89 51.46 48.24 51.55 ;
      RECT  47.51 51.96 47.96 52.1 ;
      RECT  48.69 54.48 48.98 54.77 ;
      RECT  48.68 52.87 49.5 53.04 ;
      RECT  47.95 54.62 48.24 54.77 ;
      RECT  48.75 53.98 48.92 54.48 ;
      RECT  47.79 52.1 47.96 53.75 ;
      RECT  46.98 50.54 47.33 50.89 ;
      RECT  47.09 54.48 48.24 54.62 ;
      RECT  46.68 53.57 47.25 53.9 ;
      RECT  47.89 51.55 49.51 51.72 ;
      RECT  47.51 51.78 47.68 51.96 ;
      RECT  49.22 51.49 49.51 51.55 ;
      RECT  47.45 51.49 47.74 51.78 ;
      RECT  47.73 53.98 48.02 54.04 ;
      RECT  47.73 53.75 48.02 53.81 ;
      RECT  48.96 51.19 49.25 51.27 ;
      RECT  49.21 53.04 49.5 53.1 ;
      RECT  47.09 54.46 47.96 54.48 ;
      RECT  48.68 53.04 49.03 53.13 ;
      RECT  49.21 57.31 49.5 57.25 ;
      RECT  48.96 59.14 49.25 59.08 ;
      RECT  46.53 59.08 49.61 58.93 ;
      RECT  46.98 55.35 47.33 55.0 ;
      RECT  47.73 56.31 48.92 56.14 ;
      RECT  49.22 58.4 49.51 58.34 ;
      RECT  47.09 56.22 47.25 55.66 ;
      RECT  48.68 57.34 49.03 57.25 ;
      RECT  47.89 58.4 48.24 58.31 ;
      RECT  47.89 58.66 48.24 58.57 ;
      RECT  47.51 58.16 47.96 58.02 ;
      RECT  48.69 55.64 48.98 55.35 ;
      RECT  48.68 57.25 49.5 57.08 ;
      RECT  47.95 55.5 48.24 55.35 ;
      RECT  48.75 56.14 48.92 55.64 ;
      RECT  47.79 58.02 47.96 56.37 ;
      RECT  46.98 59.58 47.33 59.23 ;
      RECT  47.09 55.64 48.24 55.5 ;
      RECT  46.68 56.55 47.25 56.22 ;
      RECT  47.89 58.57 49.51 58.4 ;
      RECT  47.51 58.34 47.68 58.16 ;
      RECT  49.22 58.63 49.51 58.57 ;
      RECT  47.45 58.63 47.74 58.34 ;
      RECT  47.73 56.14 48.02 56.08 ;
      RECT  47.73 56.37 48.02 56.31 ;
      RECT  48.96 58.93 49.25 58.85 ;
      RECT  49.21 57.08 49.5 57.02 ;
      RECT  47.09 55.66 47.96 55.64 ;
      RECT  48.68 57.08 49.03 56.99 ;
      RECT  49.21 61.51 49.5 61.57 ;
      RECT  48.96 59.68 49.25 59.74 ;
      RECT  46.53 59.74 49.61 59.89 ;
      RECT  46.98 63.47 47.33 63.82 ;
      RECT  47.73 62.51 48.92 62.68 ;
      RECT  49.22 60.42 49.51 60.48 ;
      RECT  47.09 62.6 47.25 63.16 ;
      RECT  48.68 61.48 49.03 61.57 ;
      RECT  47.89 60.42 48.24 60.51 ;
      RECT  47.89 60.16 48.24 60.25 ;
      RECT  47.51 60.66 47.96 60.8 ;
      RECT  48.69 63.18 48.98 63.47 ;
      RECT  48.68 61.57 49.5 61.74 ;
      RECT  47.95 63.32 48.24 63.47 ;
      RECT  48.75 62.68 48.92 63.18 ;
      RECT  47.79 60.8 47.96 62.45 ;
      RECT  46.98 59.24 47.33 59.59 ;
      RECT  47.09 63.18 48.24 63.32 ;
      RECT  46.68 62.27 47.25 62.6 ;
      RECT  47.89 60.25 49.51 60.42 ;
      RECT  47.51 60.48 47.68 60.66 ;
      RECT  49.22 60.19 49.51 60.25 ;
      RECT  47.45 60.19 47.74 60.48 ;
      RECT  47.73 62.68 48.02 62.74 ;
      RECT  47.73 62.45 48.02 62.51 ;
      RECT  48.96 59.89 49.25 59.97 ;
      RECT  49.21 61.74 49.5 61.8 ;
      RECT  47.09 63.16 47.96 63.18 ;
      RECT  48.68 61.74 49.03 61.83 ;
      RECT  49.21 66.01 49.5 65.95 ;
      RECT  48.96 67.84 49.25 67.78 ;
      RECT  46.53 67.78 49.61 67.63 ;
      RECT  46.98 64.05 47.33 63.7 ;
      RECT  47.73 65.01 48.92 64.84 ;
      RECT  49.22 67.1 49.51 67.04 ;
      RECT  47.09 64.92 47.25 64.36 ;
      RECT  48.68 66.04 49.03 65.95 ;
      RECT  47.89 67.1 48.24 67.01 ;
      RECT  47.89 67.36 48.24 67.27 ;
      RECT  47.51 66.86 47.96 66.72 ;
      RECT  48.69 64.34 48.98 64.05 ;
      RECT  48.68 65.95 49.5 65.78 ;
      RECT  47.95 64.2 48.24 64.05 ;
      RECT  48.75 64.84 48.92 64.34 ;
      RECT  47.79 66.72 47.96 65.07 ;
      RECT  46.98 68.28 47.33 67.93 ;
      RECT  47.09 64.34 48.24 64.2 ;
      RECT  46.68 65.25 47.25 64.92 ;
      RECT  47.89 67.27 49.51 67.1 ;
      RECT  47.51 67.04 47.68 66.86 ;
      RECT  49.22 67.33 49.51 67.27 ;
      RECT  47.45 67.33 47.74 67.04 ;
      RECT  47.73 64.84 48.02 64.78 ;
      RECT  47.73 65.07 48.02 65.01 ;
      RECT  48.96 67.63 49.25 67.55 ;
      RECT  49.21 65.78 49.5 65.72 ;
      RECT  47.09 64.36 47.96 64.34 ;
      RECT  48.68 65.78 49.03 65.69 ;
      RECT  49.21 70.21 49.5 70.27 ;
      RECT  48.96 68.38 49.25 68.44 ;
      RECT  46.53 68.44 49.61 68.59 ;
      RECT  46.98 72.17 47.33 72.52 ;
      RECT  47.73 71.21 48.92 71.38 ;
      RECT  49.22 69.12 49.51 69.18 ;
      RECT  47.09 71.3 47.25 71.86 ;
      RECT  48.68 70.18 49.03 70.27 ;
      RECT  47.89 69.12 48.24 69.21 ;
      RECT  47.89 68.86 48.24 68.95 ;
      RECT  47.51 69.36 47.96 69.5 ;
      RECT  48.69 71.88 48.98 72.17 ;
      RECT  48.68 70.27 49.5 70.44 ;
      RECT  47.95 72.02 48.24 72.17 ;
      RECT  48.75 71.38 48.92 71.88 ;
      RECT  47.79 69.5 47.96 71.15 ;
      RECT  46.98 67.94 47.33 68.29 ;
      RECT  47.09 71.88 48.24 72.02 ;
      RECT  46.68 70.97 47.25 71.3 ;
      RECT  47.89 68.95 49.51 69.12 ;
      RECT  47.51 69.18 47.68 69.36 ;
      RECT  49.22 68.89 49.51 68.95 ;
      RECT  47.45 68.89 47.74 69.18 ;
      RECT  47.73 71.38 48.02 71.44 ;
      RECT  47.73 71.15 48.02 71.21 ;
      RECT  48.96 68.59 49.25 68.67 ;
      RECT  49.21 70.44 49.5 70.5 ;
      RECT  47.09 71.86 47.96 71.88 ;
      RECT  48.68 70.44 49.03 70.53 ;
      RECT  49.21 74.71 49.5 74.65 ;
      RECT  48.96 76.54 49.25 76.48 ;
      RECT  46.53 76.48 49.61 76.33 ;
      RECT  46.98 72.75 47.33 72.4 ;
      RECT  47.73 73.71 48.92 73.54 ;
      RECT  49.22 75.8 49.51 75.74 ;
      RECT  47.09 73.62 47.25 73.06 ;
      RECT  48.68 74.74 49.03 74.65 ;
      RECT  47.89 75.8 48.24 75.71 ;
      RECT  47.89 76.06 48.24 75.97 ;
      RECT  47.51 75.56 47.96 75.42 ;
      RECT  48.69 73.04 48.98 72.75 ;
      RECT  48.68 74.65 49.5 74.48 ;
      RECT  47.95 72.9 48.24 72.75 ;
      RECT  48.75 73.54 48.92 73.04 ;
      RECT  47.79 75.42 47.96 73.77 ;
      RECT  46.98 76.98 47.33 76.63 ;
      RECT  47.09 73.04 48.24 72.9 ;
      RECT  46.68 73.95 47.25 73.62 ;
      RECT  47.89 75.97 49.51 75.8 ;
      RECT  47.51 75.74 47.68 75.56 ;
      RECT  49.22 76.03 49.51 75.97 ;
      RECT  47.45 76.03 47.74 75.74 ;
      RECT  47.73 73.54 48.02 73.48 ;
      RECT  47.73 73.77 48.02 73.71 ;
      RECT  48.96 76.33 49.25 76.25 ;
      RECT  49.21 74.48 49.5 74.42 ;
      RECT  47.09 73.06 47.96 73.04 ;
      RECT  48.68 74.48 49.03 74.39 ;
      RECT  49.21 78.91 49.5 78.97 ;
      RECT  48.96 77.08 49.25 77.14 ;
      RECT  46.53 77.14 49.61 77.29 ;
      RECT  46.98 80.87 47.33 81.22 ;
      RECT  47.73 79.91 48.92 80.08 ;
      RECT  49.22 77.82 49.51 77.88 ;
      RECT  47.09 80.0 47.25 80.56 ;
      RECT  48.68 78.88 49.03 78.97 ;
      RECT  47.89 77.82 48.24 77.91 ;
      RECT  47.89 77.56 48.24 77.65 ;
      RECT  47.51 78.06 47.96 78.2 ;
      RECT  48.69 80.58 48.98 80.87 ;
      RECT  48.68 78.97 49.5 79.14 ;
      RECT  47.95 80.72 48.24 80.87 ;
      RECT  48.75 80.08 48.92 80.58 ;
      RECT  47.79 78.2 47.96 79.85 ;
      RECT  46.98 76.64 47.33 76.99 ;
      RECT  47.09 80.58 48.24 80.72 ;
      RECT  46.68 79.67 47.25 80.0 ;
      RECT  47.89 77.65 49.51 77.82 ;
      RECT  47.51 77.88 47.68 78.06 ;
      RECT  49.22 77.59 49.51 77.65 ;
      RECT  47.45 77.59 47.74 77.88 ;
      RECT  47.73 80.08 48.02 80.14 ;
      RECT  47.73 79.85 48.02 79.91 ;
      RECT  48.96 77.29 49.25 77.37 ;
      RECT  49.21 79.14 49.5 79.2 ;
      RECT  47.09 80.56 47.96 80.58 ;
      RECT  48.68 79.14 49.03 79.23 ;
      RECT  49.21 83.41 49.5 83.35 ;
      RECT  48.96 85.24 49.25 85.18 ;
      RECT  46.53 85.18 49.61 85.03 ;
      RECT  46.98 81.45 47.33 81.1 ;
      RECT  47.73 82.41 48.92 82.24 ;
      RECT  49.22 84.5 49.51 84.44 ;
      RECT  47.09 82.32 47.25 81.76 ;
      RECT  48.68 83.44 49.03 83.35 ;
      RECT  47.89 84.5 48.24 84.41 ;
      RECT  47.89 84.76 48.24 84.67 ;
      RECT  47.51 84.26 47.96 84.12 ;
      RECT  48.69 81.74 48.98 81.45 ;
      RECT  48.68 83.35 49.5 83.18 ;
      RECT  47.95 81.6 48.24 81.45 ;
      RECT  48.75 82.24 48.92 81.74 ;
      RECT  47.79 84.12 47.96 82.47 ;
      RECT  46.98 85.68 47.33 85.33 ;
      RECT  47.09 81.74 48.24 81.6 ;
      RECT  46.68 82.65 47.25 82.32 ;
      RECT  47.89 84.67 49.51 84.5 ;
      RECT  47.51 84.44 47.68 84.26 ;
      RECT  49.22 84.73 49.51 84.67 ;
      RECT  47.45 84.73 47.74 84.44 ;
      RECT  47.73 82.24 48.02 82.18 ;
      RECT  47.73 82.47 48.02 82.41 ;
      RECT  48.96 85.03 49.25 84.95 ;
      RECT  49.21 83.18 49.5 83.12 ;
      RECT  47.09 81.76 47.96 81.74 ;
      RECT  48.68 83.18 49.03 83.09 ;
      RECT  49.21 87.61 49.5 87.67 ;
      RECT  48.96 85.78 49.25 85.84 ;
      RECT  46.53 85.84 49.61 85.99 ;
      RECT  46.98 89.57 47.33 89.92 ;
      RECT  47.73 88.61 48.92 88.78 ;
      RECT  49.22 86.52 49.51 86.58 ;
      RECT  47.09 88.7 47.25 89.26 ;
      RECT  48.68 87.58 49.03 87.67 ;
      RECT  47.89 86.52 48.24 86.61 ;
      RECT  47.89 86.26 48.24 86.35 ;
      RECT  47.51 86.76 47.96 86.9 ;
      RECT  48.69 89.28 48.98 89.57 ;
      RECT  48.68 87.67 49.5 87.84 ;
      RECT  47.95 89.42 48.24 89.57 ;
      RECT  48.75 88.78 48.92 89.28 ;
      RECT  47.79 86.9 47.96 88.55 ;
      RECT  46.98 85.34 47.33 85.69 ;
      RECT  47.09 89.28 48.24 89.42 ;
      RECT  46.68 88.37 47.25 88.7 ;
      RECT  47.89 86.35 49.51 86.52 ;
      RECT  47.51 86.58 47.68 86.76 ;
      RECT  49.22 86.29 49.51 86.35 ;
      RECT  47.45 86.29 47.74 86.58 ;
      RECT  47.73 88.78 48.02 88.84 ;
      RECT  47.73 88.55 48.02 88.61 ;
      RECT  48.96 85.99 49.25 86.07 ;
      RECT  49.21 87.84 49.5 87.9 ;
      RECT  47.09 89.26 47.96 89.28 ;
      RECT  48.68 87.84 49.03 87.93 ;
      RECT  49.21 92.11 49.5 92.05 ;
      RECT  48.96 93.94 49.25 93.88 ;
      RECT  46.53 93.88 49.61 93.73 ;
      RECT  46.98 90.15 47.33 89.8 ;
      RECT  47.73 91.11 48.92 90.94 ;
      RECT  49.22 93.2 49.51 93.14 ;
      RECT  47.09 91.02 47.25 90.46 ;
      RECT  48.68 92.14 49.03 92.05 ;
      RECT  47.89 93.2 48.24 93.11 ;
      RECT  47.89 93.46 48.24 93.37 ;
      RECT  47.51 92.96 47.96 92.82 ;
      RECT  48.69 90.44 48.98 90.15 ;
      RECT  48.68 92.05 49.5 91.88 ;
      RECT  47.95 90.3 48.24 90.15 ;
      RECT  48.75 90.94 48.92 90.44 ;
      RECT  47.79 92.82 47.96 91.17 ;
      RECT  46.98 94.38 47.33 94.03 ;
      RECT  47.09 90.44 48.24 90.3 ;
      RECT  46.68 91.35 47.25 91.02 ;
      RECT  47.89 93.37 49.51 93.2 ;
      RECT  47.51 93.14 47.68 92.96 ;
      RECT  49.22 93.43 49.51 93.37 ;
      RECT  47.45 93.43 47.74 93.14 ;
      RECT  47.73 90.94 48.02 90.88 ;
      RECT  47.73 91.17 48.02 91.11 ;
      RECT  48.96 93.73 49.25 93.65 ;
      RECT  49.21 91.88 49.5 91.82 ;
      RECT  47.09 90.46 47.96 90.44 ;
      RECT  48.68 91.88 49.03 91.79 ;
      RECT  49.21 96.31 49.5 96.37 ;
      RECT  48.96 94.48 49.25 94.54 ;
      RECT  46.53 94.54 49.61 94.69 ;
      RECT  46.98 98.27 47.33 98.62 ;
      RECT  47.73 97.31 48.92 97.48 ;
      RECT  49.22 95.22 49.51 95.28 ;
      RECT  47.09 97.4 47.25 97.96 ;
      RECT  48.68 96.28 49.03 96.37 ;
      RECT  47.89 95.22 48.24 95.31 ;
      RECT  47.89 94.96 48.24 95.05 ;
      RECT  47.51 95.46 47.96 95.6 ;
      RECT  48.69 97.98 48.98 98.27 ;
      RECT  48.68 96.37 49.5 96.54 ;
      RECT  47.95 98.12 48.24 98.27 ;
      RECT  48.75 97.48 48.92 97.98 ;
      RECT  47.79 95.6 47.96 97.25 ;
      RECT  46.98 94.04 47.33 94.39 ;
      RECT  47.09 97.98 48.24 98.12 ;
      RECT  46.68 97.07 47.25 97.4 ;
      RECT  47.89 95.05 49.51 95.22 ;
      RECT  47.51 95.28 47.68 95.46 ;
      RECT  49.22 94.99 49.51 95.05 ;
      RECT  47.45 94.99 47.74 95.28 ;
      RECT  47.73 97.48 48.02 97.54 ;
      RECT  47.73 97.25 48.02 97.31 ;
      RECT  48.96 94.69 49.25 94.77 ;
      RECT  49.21 96.54 49.5 96.6 ;
      RECT  47.09 97.96 47.96 97.98 ;
      RECT  48.68 96.54 49.03 96.63 ;
      RECT  49.21 100.81 49.5 100.75 ;
      RECT  48.96 102.64 49.25 102.58 ;
      RECT  46.53 102.58 49.61 102.43 ;
      RECT  46.98 98.85 47.33 98.5 ;
      RECT  47.73 99.81 48.92 99.64 ;
      RECT  49.22 101.9 49.51 101.84 ;
      RECT  47.09 99.72 47.25 99.16 ;
      RECT  48.68 100.84 49.03 100.75 ;
      RECT  47.89 101.9 48.24 101.81 ;
      RECT  47.89 102.16 48.24 102.07 ;
      RECT  47.51 101.66 47.96 101.52 ;
      RECT  48.69 99.14 48.98 98.85 ;
      RECT  48.68 100.75 49.5 100.58 ;
      RECT  47.95 99.0 48.24 98.85 ;
      RECT  48.75 99.64 48.92 99.14 ;
      RECT  47.79 101.52 47.96 99.87 ;
      RECT  46.98 103.08 47.33 102.73 ;
      RECT  47.09 99.14 48.24 99.0 ;
      RECT  46.68 100.05 47.25 99.72 ;
      RECT  47.89 102.07 49.51 101.9 ;
      RECT  47.51 101.84 47.68 101.66 ;
      RECT  49.22 102.13 49.51 102.07 ;
      RECT  47.45 102.13 47.74 101.84 ;
      RECT  47.73 99.64 48.02 99.58 ;
      RECT  47.73 99.87 48.02 99.81 ;
      RECT  48.96 102.43 49.25 102.35 ;
      RECT  49.21 100.58 49.5 100.52 ;
      RECT  47.09 99.16 47.96 99.14 ;
      RECT  48.68 100.58 49.03 100.49 ;
      RECT  49.21 105.01 49.5 105.07 ;
      RECT  48.96 103.18 49.25 103.24 ;
      RECT  46.53 103.24 49.61 103.39 ;
      RECT  46.98 106.97 47.33 107.32 ;
      RECT  47.73 106.01 48.92 106.18 ;
      RECT  49.22 103.92 49.51 103.98 ;
      RECT  47.09 106.1 47.25 106.66 ;
      RECT  48.68 104.98 49.03 105.07 ;
      RECT  47.89 103.92 48.24 104.01 ;
      RECT  47.89 103.66 48.24 103.75 ;
      RECT  47.51 104.16 47.96 104.3 ;
      RECT  48.69 106.68 48.98 106.97 ;
      RECT  48.68 105.07 49.5 105.24 ;
      RECT  47.95 106.82 48.24 106.97 ;
      RECT  48.75 106.18 48.92 106.68 ;
      RECT  47.79 104.3 47.96 105.95 ;
      RECT  46.98 102.74 47.33 103.09 ;
      RECT  47.09 106.68 48.24 106.82 ;
      RECT  46.68 105.77 47.25 106.1 ;
      RECT  47.89 103.75 49.51 103.92 ;
      RECT  47.51 103.98 47.68 104.16 ;
      RECT  49.22 103.69 49.51 103.75 ;
      RECT  47.45 103.69 47.74 103.98 ;
      RECT  47.73 106.18 48.02 106.24 ;
      RECT  47.73 105.95 48.02 106.01 ;
      RECT  48.96 103.39 49.25 103.47 ;
      RECT  49.21 105.24 49.5 105.3 ;
      RECT  47.09 106.66 47.96 106.68 ;
      RECT  48.68 105.24 49.03 105.33 ;
      RECT  46.53 24.94 49.61 25.09 ;
      RECT  46.53 32.83 49.61 32.98 ;
      RECT  46.53 33.64 49.61 33.79 ;
      RECT  46.53 41.53 49.61 41.68 ;
      RECT  46.53 42.34 49.61 42.49 ;
      RECT  46.53 50.23 49.61 50.38 ;
      RECT  46.53 51.04 49.61 51.19 ;
      RECT  46.53 58.93 49.61 59.08 ;
      RECT  46.53 59.74 49.61 59.89 ;
      RECT  46.53 67.63 49.61 67.78 ;
      RECT  46.53 68.44 49.61 68.59 ;
      RECT  46.53 76.33 49.61 76.48 ;
      RECT  46.53 77.14 49.61 77.29 ;
      RECT  46.53 85.03 49.61 85.18 ;
      RECT  46.53 85.84 49.61 85.99 ;
      RECT  46.53 93.73 49.61 93.88 ;
      RECT  46.53 94.54 49.61 94.69 ;
      RECT  46.53 102.43 49.61 102.58 ;
      RECT  46.53 103.24 49.61 103.39 ;
      RECT  52.29 31.21 52.58 31.15 ;
      RECT  52.04 33.04 52.33 32.98 ;
      RECT  49.61 32.98 52.69 32.83 ;
      RECT  50.06 29.25 50.41 28.9 ;
      RECT  50.81 30.21 52.0 30.04 ;
      RECT  52.3 32.3 52.59 32.24 ;
      RECT  50.17 30.12 50.33 29.56 ;
      RECT  51.76 31.24 52.11 31.15 ;
      RECT  50.97 32.3 51.32 32.21 ;
      RECT  50.97 32.56 51.32 32.47 ;
      RECT  50.59 32.06 51.04 31.92 ;
      RECT  51.77 29.54 52.06 29.25 ;
      RECT  51.76 31.15 52.58 30.98 ;
      RECT  51.03 29.4 51.32 29.25 ;
      RECT  51.83 30.04 52.0 29.54 ;
      RECT  50.87 31.92 51.04 30.27 ;
      RECT  50.06 33.48 50.41 33.13 ;
      RECT  50.17 29.54 51.32 29.4 ;
      RECT  49.76 30.45 50.33 30.12 ;
      RECT  50.97 32.47 52.59 32.3 ;
      RECT  50.59 32.24 50.76 32.06 ;
      RECT  52.3 32.53 52.59 32.47 ;
      RECT  50.53 32.53 50.82 32.24 ;
      RECT  50.81 30.04 51.1 29.98 ;
      RECT  50.81 30.27 51.1 30.21 ;
      RECT  52.04 32.83 52.33 32.75 ;
      RECT  52.29 30.98 52.58 30.92 ;
      RECT  50.17 29.56 51.04 29.54 ;
      RECT  51.76 30.98 52.11 30.89 ;
      RECT  55.37 31.21 55.66 31.15 ;
      RECT  55.12 33.04 55.41 32.98 ;
      RECT  52.69 32.98 55.77 32.83 ;
      RECT  53.14 29.25 53.49 28.9 ;
      RECT  53.89 30.21 55.08 30.04 ;
      RECT  55.38 32.3 55.67 32.24 ;
      RECT  53.25 30.12 53.41 29.56 ;
      RECT  54.84 31.24 55.19 31.15 ;
      RECT  54.05 32.3 54.4 32.21 ;
      RECT  54.05 32.56 54.4 32.47 ;
      RECT  53.67 32.06 54.12 31.92 ;
      RECT  54.85 29.54 55.14 29.25 ;
      RECT  54.84 31.15 55.66 30.98 ;
      RECT  54.11 29.4 54.4 29.25 ;
      RECT  54.91 30.04 55.08 29.54 ;
      RECT  53.95 31.92 54.12 30.27 ;
      RECT  53.14 33.48 53.49 33.13 ;
      RECT  53.25 29.54 54.4 29.4 ;
      RECT  52.84 30.45 53.41 30.12 ;
      RECT  54.05 32.47 55.67 32.3 ;
      RECT  53.67 32.24 53.84 32.06 ;
      RECT  55.38 32.53 55.67 32.47 ;
      RECT  53.61 32.53 53.9 32.24 ;
      RECT  53.89 30.04 54.18 29.98 ;
      RECT  53.89 30.27 54.18 30.21 ;
      RECT  55.12 32.83 55.41 32.75 ;
      RECT  55.37 30.98 55.66 30.92 ;
      RECT  53.25 29.56 54.12 29.54 ;
      RECT  54.84 30.98 55.19 30.89 ;
      RECT  49.61 32.98 55.77 32.83 ;
      RECT  52.29 26.71 52.58 26.77 ;
      RECT  52.04 24.88 52.33 24.94 ;
      RECT  49.61 24.94 52.69 25.09 ;
      RECT  50.06 28.67 50.41 29.02 ;
      RECT  50.81 27.71 52.0 27.88 ;
      RECT  52.3 25.62 52.59 25.68 ;
      RECT  50.17 27.8 50.33 28.36 ;
      RECT  51.76 26.68 52.11 26.77 ;
      RECT  50.97 25.62 51.32 25.71 ;
      RECT  50.97 25.36 51.32 25.45 ;
      RECT  50.59 25.86 51.04 26.0 ;
      RECT  51.77 28.38 52.06 28.67 ;
      RECT  51.76 26.77 52.58 26.94 ;
      RECT  51.03 28.52 51.32 28.67 ;
      RECT  51.83 27.88 52.0 28.38 ;
      RECT  50.87 26.0 51.04 27.65 ;
      RECT  50.06 24.44 50.41 24.79 ;
      RECT  50.17 28.38 51.32 28.52 ;
      RECT  49.76 27.47 50.33 27.8 ;
      RECT  50.97 25.45 52.59 25.62 ;
      RECT  50.59 25.68 50.76 25.86 ;
      RECT  52.3 25.39 52.59 25.45 ;
      RECT  50.53 25.39 50.82 25.68 ;
      RECT  50.81 27.88 51.1 27.94 ;
      RECT  50.81 27.65 51.1 27.71 ;
      RECT  52.04 25.09 52.33 25.17 ;
      RECT  52.29 26.94 52.58 27.0 ;
      RECT  50.17 28.36 51.04 28.38 ;
      RECT  51.76 26.94 52.11 27.03 ;
      RECT  55.37 26.71 55.66 26.77 ;
      RECT  55.12 24.88 55.41 24.94 ;
      RECT  52.69 24.94 55.77 25.09 ;
      RECT  53.14 28.67 53.49 29.02 ;
      RECT  53.89 27.71 55.08 27.88 ;
      RECT  55.38 25.62 55.67 25.68 ;
      RECT  53.25 27.8 53.41 28.36 ;
      RECT  54.84 26.68 55.19 26.77 ;
      RECT  54.05 25.62 54.4 25.71 ;
      RECT  54.05 25.36 54.4 25.45 ;
      RECT  53.67 25.86 54.12 26.0 ;
      RECT  54.85 28.38 55.14 28.67 ;
      RECT  54.84 26.77 55.66 26.94 ;
      RECT  54.11 28.52 54.4 28.67 ;
      RECT  54.91 27.88 55.08 28.38 ;
      RECT  53.95 26.0 54.12 27.65 ;
      RECT  53.14 24.44 53.49 24.79 ;
      RECT  53.25 28.38 54.4 28.52 ;
      RECT  52.84 27.47 53.41 27.8 ;
      RECT  54.05 25.45 55.67 25.62 ;
      RECT  53.67 25.68 53.84 25.86 ;
      RECT  55.38 25.39 55.67 25.45 ;
      RECT  53.61 25.39 53.9 25.68 ;
      RECT  53.89 27.88 54.18 27.94 ;
      RECT  53.89 27.65 54.18 27.71 ;
      RECT  55.12 25.09 55.41 25.17 ;
      RECT  55.37 26.94 55.66 27.0 ;
      RECT  53.25 28.36 54.12 28.38 ;
      RECT  54.84 26.94 55.19 27.03 ;
      RECT  49.61 24.94 55.77 25.09 ;
      RECT  52.29 105.01 52.58 105.07 ;
      RECT  52.04 103.18 52.33 103.24 ;
      RECT  49.61 103.24 52.69 103.39 ;
      RECT  50.06 106.97 50.41 107.32 ;
      RECT  50.81 106.01 52.0 106.18 ;
      RECT  52.3 103.92 52.59 103.98 ;
      RECT  50.17 106.1 50.33 106.66 ;
      RECT  51.76 104.98 52.11 105.07 ;
      RECT  50.97 103.92 51.32 104.01 ;
      RECT  50.97 103.66 51.32 103.75 ;
      RECT  50.59 104.16 51.04 104.3 ;
      RECT  51.77 106.68 52.06 106.97 ;
      RECT  51.76 105.07 52.58 105.24 ;
      RECT  51.03 106.82 51.32 106.97 ;
      RECT  51.83 106.18 52.0 106.68 ;
      RECT  50.87 104.3 51.04 105.95 ;
      RECT  50.06 102.74 50.41 103.09 ;
      RECT  50.17 106.68 51.32 106.82 ;
      RECT  49.76 105.77 50.33 106.1 ;
      RECT  50.97 103.75 52.59 103.92 ;
      RECT  50.59 103.98 50.76 104.16 ;
      RECT  52.3 103.69 52.59 103.75 ;
      RECT  50.53 103.69 50.82 103.98 ;
      RECT  50.81 106.18 51.1 106.24 ;
      RECT  50.81 105.95 51.1 106.01 ;
      RECT  52.04 103.39 52.33 103.47 ;
      RECT  52.29 105.24 52.58 105.3 ;
      RECT  50.17 106.66 51.04 106.68 ;
      RECT  51.76 105.24 52.11 105.33 ;
      RECT  55.37 105.01 55.66 105.07 ;
      RECT  55.12 103.18 55.41 103.24 ;
      RECT  52.69 103.24 55.77 103.39 ;
      RECT  53.14 106.97 53.49 107.32 ;
      RECT  53.89 106.01 55.08 106.18 ;
      RECT  55.38 103.92 55.67 103.98 ;
      RECT  53.25 106.1 53.41 106.66 ;
      RECT  54.84 104.98 55.19 105.07 ;
      RECT  54.05 103.92 54.4 104.01 ;
      RECT  54.05 103.66 54.4 103.75 ;
      RECT  53.67 104.16 54.12 104.3 ;
      RECT  54.85 106.68 55.14 106.97 ;
      RECT  54.84 105.07 55.66 105.24 ;
      RECT  54.11 106.82 54.4 106.97 ;
      RECT  54.91 106.18 55.08 106.68 ;
      RECT  53.95 104.3 54.12 105.95 ;
      RECT  53.14 102.74 53.49 103.09 ;
      RECT  53.25 106.68 54.4 106.82 ;
      RECT  52.84 105.77 53.41 106.1 ;
      RECT  54.05 103.75 55.67 103.92 ;
      RECT  53.67 103.98 53.84 104.16 ;
      RECT  55.38 103.69 55.67 103.75 ;
      RECT  53.61 103.69 53.9 103.98 ;
      RECT  53.89 106.18 54.18 106.24 ;
      RECT  53.89 105.95 54.18 106.01 ;
      RECT  55.12 103.39 55.41 103.47 ;
      RECT  55.37 105.24 55.66 105.3 ;
      RECT  53.25 106.66 54.12 106.68 ;
      RECT  54.84 105.24 55.19 105.33 ;
      RECT  49.61 103.24 55.77 103.39 ;
      RECT  46.13 26.71 46.42 26.77 ;
      RECT  45.88 24.88 46.17 24.94 ;
      RECT  43.45 24.94 46.53 25.09 ;
      RECT  43.9 28.67 44.25 29.02 ;
      RECT  44.65 27.71 45.84 27.88 ;
      RECT  46.14 25.62 46.43 25.68 ;
      RECT  44.01 27.8 44.17 28.36 ;
      RECT  45.6 26.68 45.95 26.77 ;
      RECT  44.81 25.62 45.16 25.71 ;
      RECT  44.81 25.36 45.16 25.45 ;
      RECT  44.43 25.86 44.88 26.0 ;
      RECT  45.61 28.38 45.9 28.67 ;
      RECT  45.6 26.77 46.42 26.94 ;
      RECT  44.87 28.52 45.16 28.67 ;
      RECT  45.67 27.88 45.84 28.38 ;
      RECT  44.71 26.0 44.88 27.65 ;
      RECT  43.9 24.44 44.25 24.79 ;
      RECT  44.01 28.38 45.16 28.52 ;
      RECT  43.6 27.47 44.17 27.8 ;
      RECT  44.81 25.45 46.43 25.62 ;
      RECT  44.43 25.68 44.6 25.86 ;
      RECT  46.14 25.39 46.43 25.45 ;
      RECT  44.37 25.39 44.66 25.68 ;
      RECT  44.65 27.88 44.94 27.94 ;
      RECT  44.65 27.65 44.94 27.71 ;
      RECT  45.88 25.09 46.17 25.17 ;
      RECT  46.13 26.94 46.42 27.0 ;
      RECT  44.01 28.36 44.88 28.38 ;
      RECT  45.6 26.94 45.95 27.03 ;
      RECT  46.13 31.21 46.42 31.15 ;
      RECT  45.88 33.04 46.17 32.98 ;
      RECT  43.45 32.98 46.53 32.83 ;
      RECT  43.9 29.25 44.25 28.9 ;
      RECT  44.65 30.21 45.84 30.04 ;
      RECT  46.14 32.3 46.43 32.24 ;
      RECT  44.01 30.12 44.17 29.56 ;
      RECT  45.6 31.24 45.95 31.15 ;
      RECT  44.81 32.3 45.16 32.21 ;
      RECT  44.81 32.56 45.16 32.47 ;
      RECT  44.43 32.06 44.88 31.92 ;
      RECT  45.61 29.54 45.9 29.25 ;
      RECT  45.6 31.15 46.42 30.98 ;
      RECT  44.87 29.4 45.16 29.25 ;
      RECT  45.67 30.04 45.84 29.54 ;
      RECT  44.71 31.92 44.88 30.27 ;
      RECT  43.9 33.48 44.25 33.13 ;
      RECT  44.01 29.54 45.16 29.4 ;
      RECT  43.6 30.45 44.17 30.12 ;
      RECT  44.81 32.47 46.43 32.3 ;
      RECT  44.43 32.24 44.6 32.06 ;
      RECT  46.14 32.53 46.43 32.47 ;
      RECT  44.37 32.53 44.66 32.24 ;
      RECT  44.65 30.04 44.94 29.98 ;
      RECT  44.65 30.27 44.94 30.21 ;
      RECT  45.88 32.83 46.17 32.75 ;
      RECT  46.13 30.98 46.42 30.92 ;
      RECT  44.01 29.56 44.88 29.54 ;
      RECT  45.6 30.98 45.95 30.89 ;
      RECT  46.13 35.41 46.42 35.47 ;
      RECT  45.88 33.58 46.17 33.64 ;
      RECT  43.45 33.64 46.53 33.79 ;
      RECT  43.9 37.37 44.25 37.72 ;
      RECT  44.65 36.41 45.84 36.58 ;
      RECT  46.14 34.32 46.43 34.38 ;
      RECT  44.01 36.5 44.17 37.06 ;
      RECT  45.6 35.38 45.95 35.47 ;
      RECT  44.81 34.32 45.16 34.41 ;
      RECT  44.81 34.06 45.16 34.15 ;
      RECT  44.43 34.56 44.88 34.7 ;
      RECT  45.61 37.08 45.9 37.37 ;
      RECT  45.6 35.47 46.42 35.64 ;
      RECT  44.87 37.22 45.16 37.37 ;
      RECT  45.67 36.58 45.84 37.08 ;
      RECT  44.71 34.7 44.88 36.35 ;
      RECT  43.9 33.14 44.25 33.49 ;
      RECT  44.01 37.08 45.16 37.22 ;
      RECT  43.6 36.17 44.17 36.5 ;
      RECT  44.81 34.15 46.43 34.32 ;
      RECT  44.43 34.38 44.6 34.56 ;
      RECT  46.14 34.09 46.43 34.15 ;
      RECT  44.37 34.09 44.66 34.38 ;
      RECT  44.65 36.58 44.94 36.64 ;
      RECT  44.65 36.35 44.94 36.41 ;
      RECT  45.88 33.79 46.17 33.87 ;
      RECT  46.13 35.64 46.42 35.7 ;
      RECT  44.01 37.06 44.88 37.08 ;
      RECT  45.6 35.64 45.95 35.73 ;
      RECT  46.13 39.91 46.42 39.85 ;
      RECT  45.88 41.74 46.17 41.68 ;
      RECT  43.45 41.68 46.53 41.53 ;
      RECT  43.9 37.95 44.25 37.6 ;
      RECT  44.65 38.91 45.84 38.74 ;
      RECT  46.14 41.0 46.43 40.94 ;
      RECT  44.01 38.82 44.17 38.26 ;
      RECT  45.6 39.94 45.95 39.85 ;
      RECT  44.81 41.0 45.16 40.91 ;
      RECT  44.81 41.26 45.16 41.17 ;
      RECT  44.43 40.76 44.88 40.62 ;
      RECT  45.61 38.24 45.9 37.95 ;
      RECT  45.6 39.85 46.42 39.68 ;
      RECT  44.87 38.1 45.16 37.95 ;
      RECT  45.67 38.74 45.84 38.24 ;
      RECT  44.71 40.62 44.88 38.97 ;
      RECT  43.9 42.18 44.25 41.83 ;
      RECT  44.01 38.24 45.16 38.1 ;
      RECT  43.6 39.15 44.17 38.82 ;
      RECT  44.81 41.17 46.43 41.0 ;
      RECT  44.43 40.94 44.6 40.76 ;
      RECT  46.14 41.23 46.43 41.17 ;
      RECT  44.37 41.23 44.66 40.94 ;
      RECT  44.65 38.74 44.94 38.68 ;
      RECT  44.65 38.97 44.94 38.91 ;
      RECT  45.88 41.53 46.17 41.45 ;
      RECT  46.13 39.68 46.42 39.62 ;
      RECT  44.01 38.26 44.88 38.24 ;
      RECT  45.6 39.68 45.95 39.59 ;
      RECT  46.13 44.11 46.42 44.17 ;
      RECT  45.88 42.28 46.17 42.34 ;
      RECT  43.45 42.34 46.53 42.49 ;
      RECT  43.9 46.07 44.25 46.42 ;
      RECT  44.65 45.11 45.84 45.28 ;
      RECT  46.14 43.02 46.43 43.08 ;
      RECT  44.01 45.2 44.17 45.76 ;
      RECT  45.6 44.08 45.95 44.17 ;
      RECT  44.81 43.02 45.16 43.11 ;
      RECT  44.81 42.76 45.16 42.85 ;
      RECT  44.43 43.26 44.88 43.4 ;
      RECT  45.61 45.78 45.9 46.07 ;
      RECT  45.6 44.17 46.42 44.34 ;
      RECT  44.87 45.92 45.16 46.07 ;
      RECT  45.67 45.28 45.84 45.78 ;
      RECT  44.71 43.4 44.88 45.05 ;
      RECT  43.9 41.84 44.25 42.19 ;
      RECT  44.01 45.78 45.16 45.92 ;
      RECT  43.6 44.87 44.17 45.2 ;
      RECT  44.81 42.85 46.43 43.02 ;
      RECT  44.43 43.08 44.6 43.26 ;
      RECT  46.14 42.79 46.43 42.85 ;
      RECT  44.37 42.79 44.66 43.08 ;
      RECT  44.65 45.28 44.94 45.34 ;
      RECT  44.65 45.05 44.94 45.11 ;
      RECT  45.88 42.49 46.17 42.57 ;
      RECT  46.13 44.34 46.42 44.4 ;
      RECT  44.01 45.76 44.88 45.78 ;
      RECT  45.6 44.34 45.95 44.43 ;
      RECT  46.13 48.61 46.42 48.55 ;
      RECT  45.88 50.44 46.17 50.38 ;
      RECT  43.45 50.38 46.53 50.23 ;
      RECT  43.9 46.65 44.25 46.3 ;
      RECT  44.65 47.61 45.84 47.44 ;
      RECT  46.14 49.7 46.43 49.64 ;
      RECT  44.01 47.52 44.17 46.96 ;
      RECT  45.6 48.64 45.95 48.55 ;
      RECT  44.81 49.7 45.16 49.61 ;
      RECT  44.81 49.96 45.16 49.87 ;
      RECT  44.43 49.46 44.88 49.32 ;
      RECT  45.61 46.94 45.9 46.65 ;
      RECT  45.6 48.55 46.42 48.38 ;
      RECT  44.87 46.8 45.16 46.65 ;
      RECT  45.67 47.44 45.84 46.94 ;
      RECT  44.71 49.32 44.88 47.67 ;
      RECT  43.9 50.88 44.25 50.53 ;
      RECT  44.01 46.94 45.16 46.8 ;
      RECT  43.6 47.85 44.17 47.52 ;
      RECT  44.81 49.87 46.43 49.7 ;
      RECT  44.43 49.64 44.6 49.46 ;
      RECT  46.14 49.93 46.43 49.87 ;
      RECT  44.37 49.93 44.66 49.64 ;
      RECT  44.65 47.44 44.94 47.38 ;
      RECT  44.65 47.67 44.94 47.61 ;
      RECT  45.88 50.23 46.17 50.15 ;
      RECT  46.13 48.38 46.42 48.32 ;
      RECT  44.01 46.96 44.88 46.94 ;
      RECT  45.6 48.38 45.95 48.29 ;
      RECT  46.13 52.81 46.42 52.87 ;
      RECT  45.88 50.98 46.17 51.04 ;
      RECT  43.45 51.04 46.53 51.19 ;
      RECT  43.9 54.77 44.25 55.12 ;
      RECT  44.65 53.81 45.84 53.98 ;
      RECT  46.14 51.72 46.43 51.78 ;
      RECT  44.01 53.9 44.17 54.46 ;
      RECT  45.6 52.78 45.95 52.87 ;
      RECT  44.81 51.72 45.16 51.81 ;
      RECT  44.81 51.46 45.16 51.55 ;
      RECT  44.43 51.96 44.88 52.1 ;
      RECT  45.61 54.48 45.9 54.77 ;
      RECT  45.6 52.87 46.42 53.04 ;
      RECT  44.87 54.62 45.16 54.77 ;
      RECT  45.67 53.98 45.84 54.48 ;
      RECT  44.71 52.1 44.88 53.75 ;
      RECT  43.9 50.54 44.25 50.89 ;
      RECT  44.01 54.48 45.16 54.62 ;
      RECT  43.6 53.57 44.17 53.9 ;
      RECT  44.81 51.55 46.43 51.72 ;
      RECT  44.43 51.78 44.6 51.96 ;
      RECT  46.14 51.49 46.43 51.55 ;
      RECT  44.37 51.49 44.66 51.78 ;
      RECT  44.65 53.98 44.94 54.04 ;
      RECT  44.65 53.75 44.94 53.81 ;
      RECT  45.88 51.19 46.17 51.27 ;
      RECT  46.13 53.04 46.42 53.1 ;
      RECT  44.01 54.46 44.88 54.48 ;
      RECT  45.6 53.04 45.95 53.13 ;
      RECT  46.13 57.31 46.42 57.25 ;
      RECT  45.88 59.14 46.17 59.08 ;
      RECT  43.45 59.08 46.53 58.93 ;
      RECT  43.9 55.35 44.25 55.0 ;
      RECT  44.65 56.31 45.84 56.14 ;
      RECT  46.14 58.4 46.43 58.34 ;
      RECT  44.01 56.22 44.17 55.66 ;
      RECT  45.6 57.34 45.95 57.25 ;
      RECT  44.81 58.4 45.16 58.31 ;
      RECT  44.81 58.66 45.16 58.57 ;
      RECT  44.43 58.16 44.88 58.02 ;
      RECT  45.61 55.64 45.9 55.35 ;
      RECT  45.6 57.25 46.42 57.08 ;
      RECT  44.87 55.5 45.16 55.35 ;
      RECT  45.67 56.14 45.84 55.64 ;
      RECT  44.71 58.02 44.88 56.37 ;
      RECT  43.9 59.58 44.25 59.23 ;
      RECT  44.01 55.64 45.16 55.5 ;
      RECT  43.6 56.55 44.17 56.22 ;
      RECT  44.81 58.57 46.43 58.4 ;
      RECT  44.43 58.34 44.6 58.16 ;
      RECT  46.14 58.63 46.43 58.57 ;
      RECT  44.37 58.63 44.66 58.34 ;
      RECT  44.65 56.14 44.94 56.08 ;
      RECT  44.65 56.37 44.94 56.31 ;
      RECT  45.88 58.93 46.17 58.85 ;
      RECT  46.13 57.08 46.42 57.02 ;
      RECT  44.01 55.66 44.88 55.64 ;
      RECT  45.6 57.08 45.95 56.99 ;
      RECT  46.13 61.51 46.42 61.57 ;
      RECT  45.88 59.68 46.17 59.74 ;
      RECT  43.45 59.74 46.53 59.89 ;
      RECT  43.9 63.47 44.25 63.82 ;
      RECT  44.65 62.51 45.84 62.68 ;
      RECT  46.14 60.42 46.43 60.48 ;
      RECT  44.01 62.6 44.17 63.16 ;
      RECT  45.6 61.48 45.95 61.57 ;
      RECT  44.81 60.42 45.16 60.51 ;
      RECT  44.81 60.16 45.16 60.25 ;
      RECT  44.43 60.66 44.88 60.8 ;
      RECT  45.61 63.18 45.9 63.47 ;
      RECT  45.6 61.57 46.42 61.74 ;
      RECT  44.87 63.32 45.16 63.47 ;
      RECT  45.67 62.68 45.84 63.18 ;
      RECT  44.71 60.8 44.88 62.45 ;
      RECT  43.9 59.24 44.25 59.59 ;
      RECT  44.01 63.18 45.16 63.32 ;
      RECT  43.6 62.27 44.17 62.6 ;
      RECT  44.81 60.25 46.43 60.42 ;
      RECT  44.43 60.48 44.6 60.66 ;
      RECT  46.14 60.19 46.43 60.25 ;
      RECT  44.37 60.19 44.66 60.48 ;
      RECT  44.65 62.68 44.94 62.74 ;
      RECT  44.65 62.45 44.94 62.51 ;
      RECT  45.88 59.89 46.17 59.97 ;
      RECT  46.13 61.74 46.42 61.8 ;
      RECT  44.01 63.16 44.88 63.18 ;
      RECT  45.6 61.74 45.95 61.83 ;
      RECT  46.13 66.01 46.42 65.95 ;
      RECT  45.88 67.84 46.17 67.78 ;
      RECT  43.45 67.78 46.53 67.63 ;
      RECT  43.9 64.05 44.25 63.7 ;
      RECT  44.65 65.01 45.84 64.84 ;
      RECT  46.14 67.1 46.43 67.04 ;
      RECT  44.01 64.92 44.17 64.36 ;
      RECT  45.6 66.04 45.95 65.95 ;
      RECT  44.81 67.1 45.16 67.01 ;
      RECT  44.81 67.36 45.16 67.27 ;
      RECT  44.43 66.86 44.88 66.72 ;
      RECT  45.61 64.34 45.9 64.05 ;
      RECT  45.6 65.95 46.42 65.78 ;
      RECT  44.87 64.2 45.16 64.05 ;
      RECT  45.67 64.84 45.84 64.34 ;
      RECT  44.71 66.72 44.88 65.07 ;
      RECT  43.9 68.28 44.25 67.93 ;
      RECT  44.01 64.34 45.16 64.2 ;
      RECT  43.6 65.25 44.17 64.92 ;
      RECT  44.81 67.27 46.43 67.1 ;
      RECT  44.43 67.04 44.6 66.86 ;
      RECT  46.14 67.33 46.43 67.27 ;
      RECT  44.37 67.33 44.66 67.04 ;
      RECT  44.65 64.84 44.94 64.78 ;
      RECT  44.65 65.07 44.94 65.01 ;
      RECT  45.88 67.63 46.17 67.55 ;
      RECT  46.13 65.78 46.42 65.72 ;
      RECT  44.01 64.36 44.88 64.34 ;
      RECT  45.6 65.78 45.95 65.69 ;
      RECT  46.13 70.21 46.42 70.27 ;
      RECT  45.88 68.38 46.17 68.44 ;
      RECT  43.45 68.44 46.53 68.59 ;
      RECT  43.9 72.17 44.25 72.52 ;
      RECT  44.65 71.21 45.84 71.38 ;
      RECT  46.14 69.12 46.43 69.18 ;
      RECT  44.01 71.3 44.17 71.86 ;
      RECT  45.6 70.18 45.95 70.27 ;
      RECT  44.81 69.12 45.16 69.21 ;
      RECT  44.81 68.86 45.16 68.95 ;
      RECT  44.43 69.36 44.88 69.5 ;
      RECT  45.61 71.88 45.9 72.17 ;
      RECT  45.6 70.27 46.42 70.44 ;
      RECT  44.87 72.02 45.16 72.17 ;
      RECT  45.67 71.38 45.84 71.88 ;
      RECT  44.71 69.5 44.88 71.15 ;
      RECT  43.9 67.94 44.25 68.29 ;
      RECT  44.01 71.88 45.16 72.02 ;
      RECT  43.6 70.97 44.17 71.3 ;
      RECT  44.81 68.95 46.43 69.12 ;
      RECT  44.43 69.18 44.6 69.36 ;
      RECT  46.14 68.89 46.43 68.95 ;
      RECT  44.37 68.89 44.66 69.18 ;
      RECT  44.65 71.38 44.94 71.44 ;
      RECT  44.65 71.15 44.94 71.21 ;
      RECT  45.88 68.59 46.17 68.67 ;
      RECT  46.13 70.44 46.42 70.5 ;
      RECT  44.01 71.86 44.88 71.88 ;
      RECT  45.6 70.44 45.95 70.53 ;
      RECT  46.13 74.71 46.42 74.65 ;
      RECT  45.88 76.54 46.17 76.48 ;
      RECT  43.45 76.48 46.53 76.33 ;
      RECT  43.9 72.75 44.25 72.4 ;
      RECT  44.65 73.71 45.84 73.54 ;
      RECT  46.14 75.8 46.43 75.74 ;
      RECT  44.01 73.62 44.17 73.06 ;
      RECT  45.6 74.74 45.95 74.65 ;
      RECT  44.81 75.8 45.16 75.71 ;
      RECT  44.81 76.06 45.16 75.97 ;
      RECT  44.43 75.56 44.88 75.42 ;
      RECT  45.61 73.04 45.9 72.75 ;
      RECT  45.6 74.65 46.42 74.48 ;
      RECT  44.87 72.9 45.16 72.75 ;
      RECT  45.67 73.54 45.84 73.04 ;
      RECT  44.71 75.42 44.88 73.77 ;
      RECT  43.9 76.98 44.25 76.63 ;
      RECT  44.01 73.04 45.16 72.9 ;
      RECT  43.6 73.95 44.17 73.62 ;
      RECT  44.81 75.97 46.43 75.8 ;
      RECT  44.43 75.74 44.6 75.56 ;
      RECT  46.14 76.03 46.43 75.97 ;
      RECT  44.37 76.03 44.66 75.74 ;
      RECT  44.65 73.54 44.94 73.48 ;
      RECT  44.65 73.77 44.94 73.71 ;
      RECT  45.88 76.33 46.17 76.25 ;
      RECT  46.13 74.48 46.42 74.42 ;
      RECT  44.01 73.06 44.88 73.04 ;
      RECT  45.6 74.48 45.95 74.39 ;
      RECT  46.13 78.91 46.42 78.97 ;
      RECT  45.88 77.08 46.17 77.14 ;
      RECT  43.45 77.14 46.53 77.29 ;
      RECT  43.9 80.87 44.25 81.22 ;
      RECT  44.65 79.91 45.84 80.08 ;
      RECT  46.14 77.82 46.43 77.88 ;
      RECT  44.01 80.0 44.17 80.56 ;
      RECT  45.6 78.88 45.95 78.97 ;
      RECT  44.81 77.82 45.16 77.91 ;
      RECT  44.81 77.56 45.16 77.65 ;
      RECT  44.43 78.06 44.88 78.2 ;
      RECT  45.61 80.58 45.9 80.87 ;
      RECT  45.6 78.97 46.42 79.14 ;
      RECT  44.87 80.72 45.16 80.87 ;
      RECT  45.67 80.08 45.84 80.58 ;
      RECT  44.71 78.2 44.88 79.85 ;
      RECT  43.9 76.64 44.25 76.99 ;
      RECT  44.01 80.58 45.16 80.72 ;
      RECT  43.6 79.67 44.17 80.0 ;
      RECT  44.81 77.65 46.43 77.82 ;
      RECT  44.43 77.88 44.6 78.06 ;
      RECT  46.14 77.59 46.43 77.65 ;
      RECT  44.37 77.59 44.66 77.88 ;
      RECT  44.65 80.08 44.94 80.14 ;
      RECT  44.65 79.85 44.94 79.91 ;
      RECT  45.88 77.29 46.17 77.37 ;
      RECT  46.13 79.14 46.42 79.2 ;
      RECT  44.01 80.56 44.88 80.58 ;
      RECT  45.6 79.14 45.95 79.23 ;
      RECT  46.13 83.41 46.42 83.35 ;
      RECT  45.88 85.24 46.17 85.18 ;
      RECT  43.45 85.18 46.53 85.03 ;
      RECT  43.9 81.45 44.25 81.1 ;
      RECT  44.65 82.41 45.84 82.24 ;
      RECT  46.14 84.5 46.43 84.44 ;
      RECT  44.01 82.32 44.17 81.76 ;
      RECT  45.6 83.44 45.95 83.35 ;
      RECT  44.81 84.5 45.16 84.41 ;
      RECT  44.81 84.76 45.16 84.67 ;
      RECT  44.43 84.26 44.88 84.12 ;
      RECT  45.61 81.74 45.9 81.45 ;
      RECT  45.6 83.35 46.42 83.18 ;
      RECT  44.87 81.6 45.16 81.45 ;
      RECT  45.67 82.24 45.84 81.74 ;
      RECT  44.71 84.12 44.88 82.47 ;
      RECT  43.9 85.68 44.25 85.33 ;
      RECT  44.01 81.74 45.16 81.6 ;
      RECT  43.6 82.65 44.17 82.32 ;
      RECT  44.81 84.67 46.43 84.5 ;
      RECT  44.43 84.44 44.6 84.26 ;
      RECT  46.14 84.73 46.43 84.67 ;
      RECT  44.37 84.73 44.66 84.44 ;
      RECT  44.65 82.24 44.94 82.18 ;
      RECT  44.65 82.47 44.94 82.41 ;
      RECT  45.88 85.03 46.17 84.95 ;
      RECT  46.13 83.18 46.42 83.12 ;
      RECT  44.01 81.76 44.88 81.74 ;
      RECT  45.6 83.18 45.95 83.09 ;
      RECT  46.13 87.61 46.42 87.67 ;
      RECT  45.88 85.78 46.17 85.84 ;
      RECT  43.45 85.84 46.53 85.99 ;
      RECT  43.9 89.57 44.25 89.92 ;
      RECT  44.65 88.61 45.84 88.78 ;
      RECT  46.14 86.52 46.43 86.58 ;
      RECT  44.01 88.7 44.17 89.26 ;
      RECT  45.6 87.58 45.95 87.67 ;
      RECT  44.81 86.52 45.16 86.61 ;
      RECT  44.81 86.26 45.16 86.35 ;
      RECT  44.43 86.76 44.88 86.9 ;
      RECT  45.61 89.28 45.9 89.57 ;
      RECT  45.6 87.67 46.42 87.84 ;
      RECT  44.87 89.42 45.16 89.57 ;
      RECT  45.67 88.78 45.84 89.28 ;
      RECT  44.71 86.9 44.88 88.55 ;
      RECT  43.9 85.34 44.25 85.69 ;
      RECT  44.01 89.28 45.16 89.42 ;
      RECT  43.6 88.37 44.17 88.7 ;
      RECT  44.81 86.35 46.43 86.52 ;
      RECT  44.43 86.58 44.6 86.76 ;
      RECT  46.14 86.29 46.43 86.35 ;
      RECT  44.37 86.29 44.66 86.58 ;
      RECT  44.65 88.78 44.94 88.84 ;
      RECT  44.65 88.55 44.94 88.61 ;
      RECT  45.88 85.99 46.17 86.07 ;
      RECT  46.13 87.84 46.42 87.9 ;
      RECT  44.01 89.26 44.88 89.28 ;
      RECT  45.6 87.84 45.95 87.93 ;
      RECT  46.13 92.11 46.42 92.05 ;
      RECT  45.88 93.94 46.17 93.88 ;
      RECT  43.45 93.88 46.53 93.73 ;
      RECT  43.9 90.15 44.25 89.8 ;
      RECT  44.65 91.11 45.84 90.94 ;
      RECT  46.14 93.2 46.43 93.14 ;
      RECT  44.01 91.02 44.17 90.46 ;
      RECT  45.6 92.14 45.95 92.05 ;
      RECT  44.81 93.2 45.16 93.11 ;
      RECT  44.81 93.46 45.16 93.37 ;
      RECT  44.43 92.96 44.88 92.82 ;
      RECT  45.61 90.44 45.9 90.15 ;
      RECT  45.6 92.05 46.42 91.88 ;
      RECT  44.87 90.3 45.16 90.15 ;
      RECT  45.67 90.94 45.84 90.44 ;
      RECT  44.71 92.82 44.88 91.17 ;
      RECT  43.9 94.38 44.25 94.03 ;
      RECT  44.01 90.44 45.16 90.3 ;
      RECT  43.6 91.35 44.17 91.02 ;
      RECT  44.81 93.37 46.43 93.2 ;
      RECT  44.43 93.14 44.6 92.96 ;
      RECT  46.14 93.43 46.43 93.37 ;
      RECT  44.37 93.43 44.66 93.14 ;
      RECT  44.65 90.94 44.94 90.88 ;
      RECT  44.65 91.17 44.94 91.11 ;
      RECT  45.88 93.73 46.17 93.65 ;
      RECT  46.13 91.88 46.42 91.82 ;
      RECT  44.01 90.46 44.88 90.44 ;
      RECT  45.6 91.88 45.95 91.79 ;
      RECT  46.13 96.31 46.42 96.37 ;
      RECT  45.88 94.48 46.17 94.54 ;
      RECT  43.45 94.54 46.53 94.69 ;
      RECT  43.9 98.27 44.25 98.62 ;
      RECT  44.65 97.31 45.84 97.48 ;
      RECT  46.14 95.22 46.43 95.28 ;
      RECT  44.01 97.4 44.17 97.96 ;
      RECT  45.6 96.28 45.95 96.37 ;
      RECT  44.81 95.22 45.16 95.31 ;
      RECT  44.81 94.96 45.16 95.05 ;
      RECT  44.43 95.46 44.88 95.6 ;
      RECT  45.61 97.98 45.9 98.27 ;
      RECT  45.6 96.37 46.42 96.54 ;
      RECT  44.87 98.12 45.16 98.27 ;
      RECT  45.67 97.48 45.84 97.98 ;
      RECT  44.71 95.6 44.88 97.25 ;
      RECT  43.9 94.04 44.25 94.39 ;
      RECT  44.01 97.98 45.16 98.12 ;
      RECT  43.6 97.07 44.17 97.4 ;
      RECT  44.81 95.05 46.43 95.22 ;
      RECT  44.43 95.28 44.6 95.46 ;
      RECT  46.14 94.99 46.43 95.05 ;
      RECT  44.37 94.99 44.66 95.28 ;
      RECT  44.65 97.48 44.94 97.54 ;
      RECT  44.65 97.25 44.94 97.31 ;
      RECT  45.88 94.69 46.17 94.77 ;
      RECT  46.13 96.54 46.42 96.6 ;
      RECT  44.01 97.96 44.88 97.98 ;
      RECT  45.6 96.54 45.95 96.63 ;
      RECT  46.13 100.81 46.42 100.75 ;
      RECT  45.88 102.64 46.17 102.58 ;
      RECT  43.45 102.58 46.53 102.43 ;
      RECT  43.9 98.85 44.25 98.5 ;
      RECT  44.65 99.81 45.84 99.64 ;
      RECT  46.14 101.9 46.43 101.84 ;
      RECT  44.01 99.72 44.17 99.16 ;
      RECT  45.6 100.84 45.95 100.75 ;
      RECT  44.81 101.9 45.16 101.81 ;
      RECT  44.81 102.16 45.16 102.07 ;
      RECT  44.43 101.66 44.88 101.52 ;
      RECT  45.61 99.14 45.9 98.85 ;
      RECT  45.6 100.75 46.42 100.58 ;
      RECT  44.87 99.0 45.16 98.85 ;
      RECT  45.67 99.64 45.84 99.14 ;
      RECT  44.71 101.52 44.88 99.87 ;
      RECT  43.9 103.08 44.25 102.73 ;
      RECT  44.01 99.14 45.16 99.0 ;
      RECT  43.6 100.05 44.17 99.72 ;
      RECT  44.81 102.07 46.43 101.9 ;
      RECT  44.43 101.84 44.6 101.66 ;
      RECT  46.14 102.13 46.43 102.07 ;
      RECT  44.37 102.13 44.66 101.84 ;
      RECT  44.65 99.64 44.94 99.58 ;
      RECT  44.65 99.87 44.94 99.81 ;
      RECT  45.88 102.43 46.17 102.35 ;
      RECT  46.13 100.58 46.42 100.52 ;
      RECT  44.01 99.16 44.88 99.14 ;
      RECT  45.6 100.58 45.95 100.49 ;
      RECT  46.13 105.01 46.42 105.07 ;
      RECT  45.88 103.18 46.17 103.24 ;
      RECT  43.45 103.24 46.53 103.39 ;
      RECT  43.9 106.97 44.25 107.32 ;
      RECT  44.65 106.01 45.84 106.18 ;
      RECT  46.14 103.92 46.43 103.98 ;
      RECT  44.01 106.1 44.17 106.66 ;
      RECT  45.6 104.98 45.95 105.07 ;
      RECT  44.81 103.92 45.16 104.01 ;
      RECT  44.81 103.66 45.16 103.75 ;
      RECT  44.43 104.16 44.88 104.3 ;
      RECT  45.61 106.68 45.9 106.97 ;
      RECT  45.6 105.07 46.42 105.24 ;
      RECT  44.87 106.82 45.16 106.97 ;
      RECT  45.67 106.18 45.84 106.68 ;
      RECT  44.71 104.3 44.88 105.95 ;
      RECT  43.9 102.74 44.25 103.09 ;
      RECT  44.01 106.68 45.16 106.82 ;
      RECT  43.6 105.77 44.17 106.1 ;
      RECT  44.81 103.75 46.43 103.92 ;
      RECT  44.43 103.98 44.6 104.16 ;
      RECT  46.14 103.69 46.43 103.75 ;
      RECT  44.37 103.69 44.66 103.98 ;
      RECT  44.65 106.18 44.94 106.24 ;
      RECT  44.65 105.95 44.94 106.01 ;
      RECT  45.88 103.39 46.17 103.47 ;
      RECT  46.13 105.24 46.42 105.3 ;
      RECT  44.01 106.66 44.88 106.68 ;
      RECT  45.6 105.24 45.95 105.33 ;
      RECT  43.45 24.94 46.53 25.09 ;
      RECT  43.45 32.83 46.53 32.98 ;
      RECT  43.45 33.64 46.53 33.79 ;
      RECT  43.45 41.53 46.53 41.68 ;
      RECT  43.45 42.34 46.53 42.49 ;
      RECT  43.45 50.23 46.53 50.38 ;
      RECT  43.45 51.04 46.53 51.19 ;
      RECT  43.45 58.93 46.53 59.08 ;
      RECT  43.45 59.74 46.53 59.89 ;
      RECT  43.45 67.63 46.53 67.78 ;
      RECT  43.45 68.44 46.53 68.59 ;
      RECT  43.45 76.33 46.53 76.48 ;
      RECT  43.45 77.14 46.53 77.29 ;
      RECT  43.45 85.03 46.53 85.18 ;
      RECT  43.45 85.84 46.53 85.99 ;
      RECT  43.45 93.73 46.53 93.88 ;
      RECT  43.45 94.54 46.53 94.69 ;
      RECT  43.45 102.43 46.53 102.58 ;
      RECT  43.45 103.24 46.53 103.39 ;
      RECT  58.45 26.71 58.74 26.77 ;
      RECT  58.2 24.88 58.49 24.94 ;
      RECT  55.77 24.94 58.85 25.09 ;
      RECT  56.22 28.67 56.57 29.02 ;
      RECT  56.97 27.71 58.16 27.88 ;
      RECT  58.46 25.62 58.75 25.68 ;
      RECT  56.33 27.8 56.49 28.36 ;
      RECT  57.92 26.68 58.27 26.77 ;
      RECT  57.13 25.62 57.48 25.71 ;
      RECT  57.13 25.36 57.48 25.45 ;
      RECT  56.75 25.86 57.2 26.0 ;
      RECT  57.93 28.38 58.22 28.67 ;
      RECT  57.92 26.77 58.74 26.94 ;
      RECT  57.19 28.52 57.48 28.67 ;
      RECT  57.99 27.88 58.16 28.38 ;
      RECT  57.03 26.0 57.2 27.65 ;
      RECT  56.22 24.44 56.57 24.79 ;
      RECT  56.33 28.38 57.48 28.52 ;
      RECT  55.92 27.47 56.49 27.8 ;
      RECT  57.13 25.45 58.75 25.62 ;
      RECT  56.75 25.68 56.92 25.86 ;
      RECT  58.46 25.39 58.75 25.45 ;
      RECT  56.69 25.39 56.98 25.68 ;
      RECT  56.97 27.88 57.26 27.94 ;
      RECT  56.97 27.65 57.26 27.71 ;
      RECT  58.2 25.09 58.49 25.17 ;
      RECT  58.45 26.94 58.74 27.0 ;
      RECT  56.33 28.36 57.2 28.38 ;
      RECT  57.92 26.94 58.27 27.03 ;
      RECT  58.45 31.21 58.74 31.15 ;
      RECT  58.2 33.04 58.49 32.98 ;
      RECT  55.77 32.98 58.85 32.83 ;
      RECT  56.22 29.25 56.57 28.9 ;
      RECT  56.97 30.21 58.16 30.04 ;
      RECT  58.46 32.3 58.75 32.24 ;
      RECT  56.33 30.12 56.49 29.56 ;
      RECT  57.92 31.24 58.27 31.15 ;
      RECT  57.13 32.3 57.48 32.21 ;
      RECT  57.13 32.56 57.48 32.47 ;
      RECT  56.75 32.06 57.2 31.92 ;
      RECT  57.93 29.54 58.22 29.25 ;
      RECT  57.92 31.15 58.74 30.98 ;
      RECT  57.19 29.4 57.48 29.25 ;
      RECT  57.99 30.04 58.16 29.54 ;
      RECT  57.03 31.92 57.2 30.27 ;
      RECT  56.22 33.48 56.57 33.13 ;
      RECT  56.33 29.54 57.48 29.4 ;
      RECT  55.92 30.45 56.49 30.12 ;
      RECT  57.13 32.47 58.75 32.3 ;
      RECT  56.75 32.24 56.92 32.06 ;
      RECT  58.46 32.53 58.75 32.47 ;
      RECT  56.69 32.53 56.98 32.24 ;
      RECT  56.97 30.04 57.26 29.98 ;
      RECT  56.97 30.27 57.26 30.21 ;
      RECT  58.2 32.83 58.49 32.75 ;
      RECT  58.45 30.98 58.74 30.92 ;
      RECT  56.33 29.56 57.2 29.54 ;
      RECT  57.92 30.98 58.27 30.89 ;
      RECT  58.45 35.41 58.74 35.47 ;
      RECT  58.2 33.58 58.49 33.64 ;
      RECT  55.77 33.64 58.85 33.79 ;
      RECT  56.22 37.37 56.57 37.72 ;
      RECT  56.97 36.41 58.16 36.58 ;
      RECT  58.46 34.32 58.75 34.38 ;
      RECT  56.33 36.5 56.49 37.06 ;
      RECT  57.92 35.38 58.27 35.47 ;
      RECT  57.13 34.32 57.48 34.41 ;
      RECT  57.13 34.06 57.48 34.15 ;
      RECT  56.75 34.56 57.2 34.7 ;
      RECT  57.93 37.08 58.22 37.37 ;
      RECT  57.92 35.47 58.74 35.64 ;
      RECT  57.19 37.22 57.48 37.37 ;
      RECT  57.99 36.58 58.16 37.08 ;
      RECT  57.03 34.7 57.2 36.35 ;
      RECT  56.22 33.14 56.57 33.49 ;
      RECT  56.33 37.08 57.48 37.22 ;
      RECT  55.92 36.17 56.49 36.5 ;
      RECT  57.13 34.15 58.75 34.32 ;
      RECT  56.75 34.38 56.92 34.56 ;
      RECT  58.46 34.09 58.75 34.15 ;
      RECT  56.69 34.09 56.98 34.38 ;
      RECT  56.97 36.58 57.26 36.64 ;
      RECT  56.97 36.35 57.26 36.41 ;
      RECT  58.2 33.79 58.49 33.87 ;
      RECT  58.45 35.64 58.74 35.7 ;
      RECT  56.33 37.06 57.2 37.08 ;
      RECT  57.92 35.64 58.27 35.73 ;
      RECT  58.45 39.91 58.74 39.85 ;
      RECT  58.2 41.74 58.49 41.68 ;
      RECT  55.77 41.68 58.85 41.53 ;
      RECT  56.22 37.95 56.57 37.6 ;
      RECT  56.97 38.91 58.16 38.74 ;
      RECT  58.46 41.0 58.75 40.94 ;
      RECT  56.33 38.82 56.49 38.26 ;
      RECT  57.92 39.94 58.27 39.85 ;
      RECT  57.13 41.0 57.48 40.91 ;
      RECT  57.13 41.26 57.48 41.17 ;
      RECT  56.75 40.76 57.2 40.62 ;
      RECT  57.93 38.24 58.22 37.95 ;
      RECT  57.92 39.85 58.74 39.68 ;
      RECT  57.19 38.1 57.48 37.95 ;
      RECT  57.99 38.74 58.16 38.24 ;
      RECT  57.03 40.62 57.2 38.97 ;
      RECT  56.22 42.18 56.57 41.83 ;
      RECT  56.33 38.24 57.48 38.1 ;
      RECT  55.92 39.15 56.49 38.82 ;
      RECT  57.13 41.17 58.75 41.0 ;
      RECT  56.75 40.94 56.92 40.76 ;
      RECT  58.46 41.23 58.75 41.17 ;
      RECT  56.69 41.23 56.98 40.94 ;
      RECT  56.97 38.74 57.26 38.68 ;
      RECT  56.97 38.97 57.26 38.91 ;
      RECT  58.2 41.53 58.49 41.45 ;
      RECT  58.45 39.68 58.74 39.62 ;
      RECT  56.33 38.26 57.2 38.24 ;
      RECT  57.92 39.68 58.27 39.59 ;
      RECT  58.45 44.11 58.74 44.17 ;
      RECT  58.2 42.28 58.49 42.34 ;
      RECT  55.77 42.34 58.85 42.49 ;
      RECT  56.22 46.07 56.57 46.42 ;
      RECT  56.97 45.11 58.16 45.28 ;
      RECT  58.46 43.02 58.75 43.08 ;
      RECT  56.33 45.2 56.49 45.76 ;
      RECT  57.92 44.08 58.27 44.17 ;
      RECT  57.13 43.02 57.48 43.11 ;
      RECT  57.13 42.76 57.48 42.85 ;
      RECT  56.75 43.26 57.2 43.4 ;
      RECT  57.93 45.78 58.22 46.07 ;
      RECT  57.92 44.17 58.74 44.34 ;
      RECT  57.19 45.92 57.48 46.07 ;
      RECT  57.99 45.28 58.16 45.78 ;
      RECT  57.03 43.4 57.2 45.05 ;
      RECT  56.22 41.84 56.57 42.19 ;
      RECT  56.33 45.78 57.48 45.92 ;
      RECT  55.92 44.87 56.49 45.2 ;
      RECT  57.13 42.85 58.75 43.02 ;
      RECT  56.75 43.08 56.92 43.26 ;
      RECT  58.46 42.79 58.75 42.85 ;
      RECT  56.69 42.79 56.98 43.08 ;
      RECT  56.97 45.28 57.26 45.34 ;
      RECT  56.97 45.05 57.26 45.11 ;
      RECT  58.2 42.49 58.49 42.57 ;
      RECT  58.45 44.34 58.74 44.4 ;
      RECT  56.33 45.76 57.2 45.78 ;
      RECT  57.92 44.34 58.27 44.43 ;
      RECT  58.45 48.61 58.74 48.55 ;
      RECT  58.2 50.44 58.49 50.38 ;
      RECT  55.77 50.38 58.85 50.23 ;
      RECT  56.22 46.65 56.57 46.3 ;
      RECT  56.97 47.61 58.16 47.44 ;
      RECT  58.46 49.7 58.75 49.64 ;
      RECT  56.33 47.52 56.49 46.96 ;
      RECT  57.92 48.64 58.27 48.55 ;
      RECT  57.13 49.7 57.48 49.61 ;
      RECT  57.13 49.96 57.48 49.87 ;
      RECT  56.75 49.46 57.2 49.32 ;
      RECT  57.93 46.94 58.22 46.65 ;
      RECT  57.92 48.55 58.74 48.38 ;
      RECT  57.19 46.8 57.48 46.65 ;
      RECT  57.99 47.44 58.16 46.94 ;
      RECT  57.03 49.32 57.2 47.67 ;
      RECT  56.22 50.88 56.57 50.53 ;
      RECT  56.33 46.94 57.48 46.8 ;
      RECT  55.92 47.85 56.49 47.52 ;
      RECT  57.13 49.87 58.75 49.7 ;
      RECT  56.75 49.64 56.92 49.46 ;
      RECT  58.46 49.93 58.75 49.87 ;
      RECT  56.69 49.93 56.98 49.64 ;
      RECT  56.97 47.44 57.26 47.38 ;
      RECT  56.97 47.67 57.26 47.61 ;
      RECT  58.2 50.23 58.49 50.15 ;
      RECT  58.45 48.38 58.74 48.32 ;
      RECT  56.33 46.96 57.2 46.94 ;
      RECT  57.92 48.38 58.27 48.29 ;
      RECT  58.45 52.81 58.74 52.87 ;
      RECT  58.2 50.98 58.49 51.04 ;
      RECT  55.77 51.04 58.85 51.19 ;
      RECT  56.22 54.77 56.57 55.12 ;
      RECT  56.97 53.81 58.16 53.98 ;
      RECT  58.46 51.72 58.75 51.78 ;
      RECT  56.33 53.9 56.49 54.46 ;
      RECT  57.92 52.78 58.27 52.87 ;
      RECT  57.13 51.72 57.48 51.81 ;
      RECT  57.13 51.46 57.48 51.55 ;
      RECT  56.75 51.96 57.2 52.1 ;
      RECT  57.93 54.48 58.22 54.77 ;
      RECT  57.92 52.87 58.74 53.04 ;
      RECT  57.19 54.62 57.48 54.77 ;
      RECT  57.99 53.98 58.16 54.48 ;
      RECT  57.03 52.1 57.2 53.75 ;
      RECT  56.22 50.54 56.57 50.89 ;
      RECT  56.33 54.48 57.48 54.62 ;
      RECT  55.92 53.57 56.49 53.9 ;
      RECT  57.13 51.55 58.75 51.72 ;
      RECT  56.75 51.78 56.92 51.96 ;
      RECT  58.46 51.49 58.75 51.55 ;
      RECT  56.69 51.49 56.98 51.78 ;
      RECT  56.97 53.98 57.26 54.04 ;
      RECT  56.97 53.75 57.26 53.81 ;
      RECT  58.2 51.19 58.49 51.27 ;
      RECT  58.45 53.04 58.74 53.1 ;
      RECT  56.33 54.46 57.2 54.48 ;
      RECT  57.92 53.04 58.27 53.13 ;
      RECT  58.45 57.31 58.74 57.25 ;
      RECT  58.2 59.14 58.49 59.08 ;
      RECT  55.77 59.08 58.85 58.93 ;
      RECT  56.22 55.35 56.57 55.0 ;
      RECT  56.97 56.31 58.16 56.14 ;
      RECT  58.46 58.4 58.75 58.34 ;
      RECT  56.33 56.22 56.49 55.66 ;
      RECT  57.92 57.34 58.27 57.25 ;
      RECT  57.13 58.4 57.48 58.31 ;
      RECT  57.13 58.66 57.48 58.57 ;
      RECT  56.75 58.16 57.2 58.02 ;
      RECT  57.93 55.64 58.22 55.35 ;
      RECT  57.92 57.25 58.74 57.08 ;
      RECT  57.19 55.5 57.48 55.35 ;
      RECT  57.99 56.14 58.16 55.64 ;
      RECT  57.03 58.02 57.2 56.37 ;
      RECT  56.22 59.58 56.57 59.23 ;
      RECT  56.33 55.64 57.48 55.5 ;
      RECT  55.92 56.55 56.49 56.22 ;
      RECT  57.13 58.57 58.75 58.4 ;
      RECT  56.75 58.34 56.92 58.16 ;
      RECT  58.46 58.63 58.75 58.57 ;
      RECT  56.69 58.63 56.98 58.34 ;
      RECT  56.97 56.14 57.26 56.08 ;
      RECT  56.97 56.37 57.26 56.31 ;
      RECT  58.2 58.93 58.49 58.85 ;
      RECT  58.45 57.08 58.74 57.02 ;
      RECT  56.33 55.66 57.2 55.64 ;
      RECT  57.92 57.08 58.27 56.99 ;
      RECT  58.45 61.51 58.74 61.57 ;
      RECT  58.2 59.68 58.49 59.74 ;
      RECT  55.77 59.74 58.85 59.89 ;
      RECT  56.22 63.47 56.57 63.82 ;
      RECT  56.97 62.51 58.16 62.68 ;
      RECT  58.46 60.42 58.75 60.48 ;
      RECT  56.33 62.6 56.49 63.16 ;
      RECT  57.92 61.48 58.27 61.57 ;
      RECT  57.13 60.42 57.48 60.51 ;
      RECT  57.13 60.16 57.48 60.25 ;
      RECT  56.75 60.66 57.2 60.8 ;
      RECT  57.93 63.18 58.22 63.47 ;
      RECT  57.92 61.57 58.74 61.74 ;
      RECT  57.19 63.32 57.48 63.47 ;
      RECT  57.99 62.68 58.16 63.18 ;
      RECT  57.03 60.8 57.2 62.45 ;
      RECT  56.22 59.24 56.57 59.59 ;
      RECT  56.33 63.18 57.48 63.32 ;
      RECT  55.92 62.27 56.49 62.6 ;
      RECT  57.13 60.25 58.75 60.42 ;
      RECT  56.75 60.48 56.92 60.66 ;
      RECT  58.46 60.19 58.75 60.25 ;
      RECT  56.69 60.19 56.98 60.48 ;
      RECT  56.97 62.68 57.26 62.74 ;
      RECT  56.97 62.45 57.26 62.51 ;
      RECT  58.2 59.89 58.49 59.97 ;
      RECT  58.45 61.74 58.74 61.8 ;
      RECT  56.33 63.16 57.2 63.18 ;
      RECT  57.92 61.74 58.27 61.83 ;
      RECT  58.45 66.01 58.74 65.95 ;
      RECT  58.2 67.84 58.49 67.78 ;
      RECT  55.77 67.78 58.85 67.63 ;
      RECT  56.22 64.05 56.57 63.7 ;
      RECT  56.97 65.01 58.16 64.84 ;
      RECT  58.46 67.1 58.75 67.04 ;
      RECT  56.33 64.92 56.49 64.36 ;
      RECT  57.92 66.04 58.27 65.95 ;
      RECT  57.13 67.1 57.48 67.01 ;
      RECT  57.13 67.36 57.48 67.27 ;
      RECT  56.75 66.86 57.2 66.72 ;
      RECT  57.93 64.34 58.22 64.05 ;
      RECT  57.92 65.95 58.74 65.78 ;
      RECT  57.19 64.2 57.48 64.05 ;
      RECT  57.99 64.84 58.16 64.34 ;
      RECT  57.03 66.72 57.2 65.07 ;
      RECT  56.22 68.28 56.57 67.93 ;
      RECT  56.33 64.34 57.48 64.2 ;
      RECT  55.92 65.25 56.49 64.92 ;
      RECT  57.13 67.27 58.75 67.1 ;
      RECT  56.75 67.04 56.92 66.86 ;
      RECT  58.46 67.33 58.75 67.27 ;
      RECT  56.69 67.33 56.98 67.04 ;
      RECT  56.97 64.84 57.26 64.78 ;
      RECT  56.97 65.07 57.26 65.01 ;
      RECT  58.2 67.63 58.49 67.55 ;
      RECT  58.45 65.78 58.74 65.72 ;
      RECT  56.33 64.36 57.2 64.34 ;
      RECT  57.92 65.78 58.27 65.69 ;
      RECT  58.45 70.21 58.74 70.27 ;
      RECT  58.2 68.38 58.49 68.44 ;
      RECT  55.77 68.44 58.85 68.59 ;
      RECT  56.22 72.17 56.57 72.52 ;
      RECT  56.97 71.21 58.16 71.38 ;
      RECT  58.46 69.12 58.75 69.18 ;
      RECT  56.33 71.3 56.49 71.86 ;
      RECT  57.92 70.18 58.27 70.27 ;
      RECT  57.13 69.12 57.48 69.21 ;
      RECT  57.13 68.86 57.48 68.95 ;
      RECT  56.75 69.36 57.2 69.5 ;
      RECT  57.93 71.88 58.22 72.17 ;
      RECT  57.92 70.27 58.74 70.44 ;
      RECT  57.19 72.02 57.48 72.17 ;
      RECT  57.99 71.38 58.16 71.88 ;
      RECT  57.03 69.5 57.2 71.15 ;
      RECT  56.22 67.94 56.57 68.29 ;
      RECT  56.33 71.88 57.48 72.02 ;
      RECT  55.92 70.97 56.49 71.3 ;
      RECT  57.13 68.95 58.75 69.12 ;
      RECT  56.75 69.18 56.92 69.36 ;
      RECT  58.46 68.89 58.75 68.95 ;
      RECT  56.69 68.89 56.98 69.18 ;
      RECT  56.97 71.38 57.26 71.44 ;
      RECT  56.97 71.15 57.26 71.21 ;
      RECT  58.2 68.59 58.49 68.67 ;
      RECT  58.45 70.44 58.74 70.5 ;
      RECT  56.33 71.86 57.2 71.88 ;
      RECT  57.92 70.44 58.27 70.53 ;
      RECT  58.45 74.71 58.74 74.65 ;
      RECT  58.2 76.54 58.49 76.48 ;
      RECT  55.77 76.48 58.85 76.33 ;
      RECT  56.22 72.75 56.57 72.4 ;
      RECT  56.97 73.71 58.16 73.54 ;
      RECT  58.46 75.8 58.75 75.74 ;
      RECT  56.33 73.62 56.49 73.06 ;
      RECT  57.92 74.74 58.27 74.65 ;
      RECT  57.13 75.8 57.48 75.71 ;
      RECT  57.13 76.06 57.48 75.97 ;
      RECT  56.75 75.56 57.2 75.42 ;
      RECT  57.93 73.04 58.22 72.75 ;
      RECT  57.92 74.65 58.74 74.48 ;
      RECT  57.19 72.9 57.48 72.75 ;
      RECT  57.99 73.54 58.16 73.04 ;
      RECT  57.03 75.42 57.2 73.77 ;
      RECT  56.22 76.98 56.57 76.63 ;
      RECT  56.33 73.04 57.48 72.9 ;
      RECT  55.92 73.95 56.49 73.62 ;
      RECT  57.13 75.97 58.75 75.8 ;
      RECT  56.75 75.74 56.92 75.56 ;
      RECT  58.46 76.03 58.75 75.97 ;
      RECT  56.69 76.03 56.98 75.74 ;
      RECT  56.97 73.54 57.26 73.48 ;
      RECT  56.97 73.77 57.26 73.71 ;
      RECT  58.2 76.33 58.49 76.25 ;
      RECT  58.45 74.48 58.74 74.42 ;
      RECT  56.33 73.06 57.2 73.04 ;
      RECT  57.92 74.48 58.27 74.39 ;
      RECT  58.45 78.91 58.74 78.97 ;
      RECT  58.2 77.08 58.49 77.14 ;
      RECT  55.77 77.14 58.85 77.29 ;
      RECT  56.22 80.87 56.57 81.22 ;
      RECT  56.97 79.91 58.16 80.08 ;
      RECT  58.46 77.82 58.75 77.88 ;
      RECT  56.33 80.0 56.49 80.56 ;
      RECT  57.92 78.88 58.27 78.97 ;
      RECT  57.13 77.82 57.48 77.91 ;
      RECT  57.13 77.56 57.48 77.65 ;
      RECT  56.75 78.06 57.2 78.2 ;
      RECT  57.93 80.58 58.22 80.87 ;
      RECT  57.92 78.97 58.74 79.14 ;
      RECT  57.19 80.72 57.48 80.87 ;
      RECT  57.99 80.08 58.16 80.58 ;
      RECT  57.03 78.2 57.2 79.85 ;
      RECT  56.22 76.64 56.57 76.99 ;
      RECT  56.33 80.58 57.48 80.72 ;
      RECT  55.92 79.67 56.49 80.0 ;
      RECT  57.13 77.65 58.75 77.82 ;
      RECT  56.75 77.88 56.92 78.06 ;
      RECT  58.46 77.59 58.75 77.65 ;
      RECT  56.69 77.59 56.98 77.88 ;
      RECT  56.97 80.08 57.26 80.14 ;
      RECT  56.97 79.85 57.26 79.91 ;
      RECT  58.2 77.29 58.49 77.37 ;
      RECT  58.45 79.14 58.74 79.2 ;
      RECT  56.33 80.56 57.2 80.58 ;
      RECT  57.92 79.14 58.27 79.23 ;
      RECT  58.45 83.41 58.74 83.35 ;
      RECT  58.2 85.24 58.49 85.18 ;
      RECT  55.77 85.18 58.85 85.03 ;
      RECT  56.22 81.45 56.57 81.1 ;
      RECT  56.97 82.41 58.16 82.24 ;
      RECT  58.46 84.5 58.75 84.44 ;
      RECT  56.33 82.32 56.49 81.76 ;
      RECT  57.92 83.44 58.27 83.35 ;
      RECT  57.13 84.5 57.48 84.41 ;
      RECT  57.13 84.76 57.48 84.67 ;
      RECT  56.75 84.26 57.2 84.12 ;
      RECT  57.93 81.74 58.22 81.45 ;
      RECT  57.92 83.35 58.74 83.18 ;
      RECT  57.19 81.6 57.48 81.45 ;
      RECT  57.99 82.24 58.16 81.74 ;
      RECT  57.03 84.12 57.2 82.47 ;
      RECT  56.22 85.68 56.57 85.33 ;
      RECT  56.33 81.74 57.48 81.6 ;
      RECT  55.92 82.65 56.49 82.32 ;
      RECT  57.13 84.67 58.75 84.5 ;
      RECT  56.75 84.44 56.92 84.26 ;
      RECT  58.46 84.73 58.75 84.67 ;
      RECT  56.69 84.73 56.98 84.44 ;
      RECT  56.97 82.24 57.26 82.18 ;
      RECT  56.97 82.47 57.26 82.41 ;
      RECT  58.2 85.03 58.49 84.95 ;
      RECT  58.45 83.18 58.74 83.12 ;
      RECT  56.33 81.76 57.2 81.74 ;
      RECT  57.92 83.18 58.27 83.09 ;
      RECT  58.45 87.61 58.74 87.67 ;
      RECT  58.2 85.78 58.49 85.84 ;
      RECT  55.77 85.84 58.85 85.99 ;
      RECT  56.22 89.57 56.57 89.92 ;
      RECT  56.97 88.61 58.16 88.78 ;
      RECT  58.46 86.52 58.75 86.58 ;
      RECT  56.33 88.7 56.49 89.26 ;
      RECT  57.92 87.58 58.27 87.67 ;
      RECT  57.13 86.52 57.48 86.61 ;
      RECT  57.13 86.26 57.48 86.35 ;
      RECT  56.75 86.76 57.2 86.9 ;
      RECT  57.93 89.28 58.22 89.57 ;
      RECT  57.92 87.67 58.74 87.84 ;
      RECT  57.19 89.42 57.48 89.57 ;
      RECT  57.99 88.78 58.16 89.28 ;
      RECT  57.03 86.9 57.2 88.55 ;
      RECT  56.22 85.34 56.57 85.69 ;
      RECT  56.33 89.28 57.48 89.42 ;
      RECT  55.92 88.37 56.49 88.7 ;
      RECT  57.13 86.35 58.75 86.52 ;
      RECT  56.75 86.58 56.92 86.76 ;
      RECT  58.46 86.29 58.75 86.35 ;
      RECT  56.69 86.29 56.98 86.58 ;
      RECT  56.97 88.78 57.26 88.84 ;
      RECT  56.97 88.55 57.26 88.61 ;
      RECT  58.2 85.99 58.49 86.07 ;
      RECT  58.45 87.84 58.74 87.9 ;
      RECT  56.33 89.26 57.2 89.28 ;
      RECT  57.92 87.84 58.27 87.93 ;
      RECT  58.45 92.11 58.74 92.05 ;
      RECT  58.2 93.94 58.49 93.88 ;
      RECT  55.77 93.88 58.85 93.73 ;
      RECT  56.22 90.15 56.57 89.8 ;
      RECT  56.97 91.11 58.16 90.94 ;
      RECT  58.46 93.2 58.75 93.14 ;
      RECT  56.33 91.02 56.49 90.46 ;
      RECT  57.92 92.14 58.27 92.05 ;
      RECT  57.13 93.2 57.48 93.11 ;
      RECT  57.13 93.46 57.48 93.37 ;
      RECT  56.75 92.96 57.2 92.82 ;
      RECT  57.93 90.44 58.22 90.15 ;
      RECT  57.92 92.05 58.74 91.88 ;
      RECT  57.19 90.3 57.48 90.15 ;
      RECT  57.99 90.94 58.16 90.44 ;
      RECT  57.03 92.82 57.2 91.17 ;
      RECT  56.22 94.38 56.57 94.03 ;
      RECT  56.33 90.44 57.48 90.3 ;
      RECT  55.92 91.35 56.49 91.02 ;
      RECT  57.13 93.37 58.75 93.2 ;
      RECT  56.75 93.14 56.92 92.96 ;
      RECT  58.46 93.43 58.75 93.37 ;
      RECT  56.69 93.43 56.98 93.14 ;
      RECT  56.97 90.94 57.26 90.88 ;
      RECT  56.97 91.17 57.26 91.11 ;
      RECT  58.2 93.73 58.49 93.65 ;
      RECT  58.45 91.88 58.74 91.82 ;
      RECT  56.33 90.46 57.2 90.44 ;
      RECT  57.92 91.88 58.27 91.79 ;
      RECT  58.45 96.31 58.74 96.37 ;
      RECT  58.2 94.48 58.49 94.54 ;
      RECT  55.77 94.54 58.85 94.69 ;
      RECT  56.22 98.27 56.57 98.62 ;
      RECT  56.97 97.31 58.16 97.48 ;
      RECT  58.46 95.22 58.75 95.28 ;
      RECT  56.33 97.4 56.49 97.96 ;
      RECT  57.92 96.28 58.27 96.37 ;
      RECT  57.13 95.22 57.48 95.31 ;
      RECT  57.13 94.96 57.48 95.05 ;
      RECT  56.75 95.46 57.2 95.6 ;
      RECT  57.93 97.98 58.22 98.27 ;
      RECT  57.92 96.37 58.74 96.54 ;
      RECT  57.19 98.12 57.48 98.27 ;
      RECT  57.99 97.48 58.16 97.98 ;
      RECT  57.03 95.6 57.2 97.25 ;
      RECT  56.22 94.04 56.57 94.39 ;
      RECT  56.33 97.98 57.48 98.12 ;
      RECT  55.92 97.07 56.49 97.4 ;
      RECT  57.13 95.05 58.75 95.22 ;
      RECT  56.75 95.28 56.92 95.46 ;
      RECT  58.46 94.99 58.75 95.05 ;
      RECT  56.69 94.99 56.98 95.28 ;
      RECT  56.97 97.48 57.26 97.54 ;
      RECT  56.97 97.25 57.26 97.31 ;
      RECT  58.2 94.69 58.49 94.77 ;
      RECT  58.45 96.54 58.74 96.6 ;
      RECT  56.33 97.96 57.2 97.98 ;
      RECT  57.92 96.54 58.27 96.63 ;
      RECT  58.45 100.81 58.74 100.75 ;
      RECT  58.2 102.64 58.49 102.58 ;
      RECT  55.77 102.58 58.85 102.43 ;
      RECT  56.22 98.85 56.57 98.5 ;
      RECT  56.97 99.81 58.16 99.64 ;
      RECT  58.46 101.9 58.75 101.84 ;
      RECT  56.33 99.72 56.49 99.16 ;
      RECT  57.92 100.84 58.27 100.75 ;
      RECT  57.13 101.9 57.48 101.81 ;
      RECT  57.13 102.16 57.48 102.07 ;
      RECT  56.75 101.66 57.2 101.52 ;
      RECT  57.93 99.14 58.22 98.85 ;
      RECT  57.92 100.75 58.74 100.58 ;
      RECT  57.19 99.0 57.48 98.85 ;
      RECT  57.99 99.64 58.16 99.14 ;
      RECT  57.03 101.52 57.2 99.87 ;
      RECT  56.22 103.08 56.57 102.73 ;
      RECT  56.33 99.14 57.48 99.0 ;
      RECT  55.92 100.05 56.49 99.72 ;
      RECT  57.13 102.07 58.75 101.9 ;
      RECT  56.75 101.84 56.92 101.66 ;
      RECT  58.46 102.13 58.75 102.07 ;
      RECT  56.69 102.13 56.98 101.84 ;
      RECT  56.97 99.64 57.26 99.58 ;
      RECT  56.97 99.87 57.26 99.81 ;
      RECT  58.2 102.43 58.49 102.35 ;
      RECT  58.45 100.58 58.74 100.52 ;
      RECT  56.33 99.16 57.2 99.14 ;
      RECT  57.92 100.58 58.27 100.49 ;
      RECT  58.45 105.01 58.74 105.07 ;
      RECT  58.2 103.18 58.49 103.24 ;
      RECT  55.77 103.24 58.85 103.39 ;
      RECT  56.22 106.97 56.57 107.32 ;
      RECT  56.97 106.01 58.16 106.18 ;
      RECT  58.46 103.92 58.75 103.98 ;
      RECT  56.33 106.1 56.49 106.66 ;
      RECT  57.92 104.98 58.27 105.07 ;
      RECT  57.13 103.92 57.48 104.01 ;
      RECT  57.13 103.66 57.48 103.75 ;
      RECT  56.75 104.16 57.2 104.3 ;
      RECT  57.93 106.68 58.22 106.97 ;
      RECT  57.92 105.07 58.74 105.24 ;
      RECT  57.19 106.82 57.48 106.97 ;
      RECT  57.99 106.18 58.16 106.68 ;
      RECT  57.03 104.3 57.2 105.95 ;
      RECT  56.22 102.74 56.57 103.09 ;
      RECT  56.33 106.68 57.48 106.82 ;
      RECT  55.92 105.77 56.49 106.1 ;
      RECT  57.13 103.75 58.75 103.92 ;
      RECT  56.75 103.98 56.92 104.16 ;
      RECT  58.46 103.69 58.75 103.75 ;
      RECT  56.69 103.69 56.98 103.98 ;
      RECT  56.97 106.18 57.26 106.24 ;
      RECT  56.97 105.95 57.26 106.01 ;
      RECT  58.2 103.39 58.49 103.47 ;
      RECT  58.45 105.24 58.74 105.3 ;
      RECT  56.33 106.66 57.2 106.68 ;
      RECT  57.92 105.24 58.27 105.33 ;
      RECT  55.77 24.94 58.85 25.09 ;
      RECT  55.77 32.83 58.85 32.98 ;
      RECT  55.77 33.64 58.85 33.79 ;
      RECT  55.77 41.53 58.85 41.68 ;
      RECT  55.77 42.34 58.85 42.49 ;
      RECT  55.77 50.23 58.85 50.38 ;
      RECT  55.77 51.04 58.85 51.19 ;
      RECT  55.77 58.93 58.85 59.08 ;
      RECT  55.77 59.74 58.85 59.89 ;
      RECT  55.77 67.63 58.85 67.78 ;
      RECT  55.77 68.44 58.85 68.59 ;
      RECT  55.77 76.33 58.85 76.48 ;
      RECT  55.77 77.14 58.85 77.29 ;
      RECT  55.77 85.03 58.85 85.18 ;
      RECT  55.77 85.84 58.85 85.99 ;
      RECT  55.77 93.73 58.85 93.88 ;
      RECT  55.77 94.54 58.85 94.69 ;
      RECT  55.77 102.43 58.85 102.58 ;
      RECT  55.77 103.24 58.85 103.39 ;
      RECT  42.55 32.83 59.75 32.98 ;
      RECT  42.55 33.64 59.75 33.79 ;
      RECT  42.55 41.53 59.75 41.68 ;
      RECT  42.55 42.34 59.75 42.49 ;
      RECT  42.55 50.23 59.75 50.38 ;
      RECT  42.55 51.04 59.75 51.19 ;
      RECT  42.55 58.93 59.75 59.08 ;
      RECT  42.55 59.74 59.75 59.89 ;
      RECT  42.55 67.63 59.75 67.78 ;
      RECT  42.55 68.44 59.75 68.59 ;
      RECT  42.55 76.33 59.75 76.48 ;
      RECT  42.55 77.14 59.75 77.29 ;
      RECT  42.55 85.03 59.75 85.18 ;
      RECT  42.55 85.84 59.75 85.99 ;
      RECT  42.55 93.73 59.75 93.88 ;
      RECT  42.55 94.54 59.75 94.69 ;
      RECT  42.55 102.43 59.75 102.58 ;
      RECT  46.53 16.785 49.61 16.925 ;
      RECT  49.61 16.785 52.69 16.925 ;
      RECT  52.69 16.785 55.77 16.925 ;
      RECT  42.55 16.785 55.77 16.925 ;
      RECT  49.61 13.5 52.69 13.79 ;
      RECT  51.57 13.06 51.86 13.35 ;
      RECT  51.7 11.22 51.99 11.51 ;
      RECT  50.62 12.35 51.71 12.53 ;
      RECT  51.7 9.78 51.99 10.07 ;
      RECT  49.76 10.3 51.64 10.44 ;
      RECT  49.76 10.01 50.07 10.3 ;
      RECT  51.35 10.44 51.64 10.59 ;
      RECT  49.61 8.91 52.69 9.2 ;
      RECT  49.75 11.71 50.03 11.73 ;
      RECT  50.86 10.61 51.21 10.96 ;
      RECT  52.2 11.02 52.55 11.37 ;
      RECT  50.89 9.64 51.18 9.7 ;
      RECT  50.47 12.26 50.78 12.33 ;
      RECT  49.61 11.73 52.69 11.9 ;
      RECT  52.01 12.84 52.21 13.5 ;
      RECT  50.87 9.39 51.2 9.47 ;
      RECT  51.81 10.07 51.96 11.22 ;
      RECT  51.92 12.55 52.21 12.84 ;
      RECT  51.57 12.53 51.71 13.06 ;
      RECT  50.47 12.04 50.76 12.26 ;
      RECT  49.75 11.9 50.03 12.0 ;
      RECT  49.61 9.47 52.69 9.64 ;
      RECT  50.61 12.33 50.78 12.35 ;
      RECT  49.76 10.44 50.07 10.73 ;
      RECT  52.69 13.5 55.77 13.79 ;
      RECT  54.65 13.06 54.94 13.35 ;
      RECT  54.78 11.22 55.07 11.51 ;
      RECT  53.7 12.35 54.79 12.53 ;
      RECT  54.78 9.78 55.07 10.07 ;
      RECT  52.84 10.3 54.72 10.44 ;
      RECT  52.84 10.01 53.15 10.3 ;
      RECT  54.43 10.44 54.72 10.59 ;
      RECT  52.69 8.91 55.77 9.2 ;
      RECT  52.83 11.71 53.11 11.73 ;
      RECT  53.94 10.61 54.29 10.96 ;
      RECT  55.28 11.02 55.63 11.37 ;
      RECT  53.97 9.64 54.26 9.7 ;
      RECT  53.55 12.26 53.86 12.33 ;
      RECT  52.69 11.73 55.77 11.9 ;
      RECT  55.09 12.84 55.29 13.5 ;
      RECT  53.95 9.39 54.28 9.47 ;
      RECT  54.89 10.07 55.04 11.22 ;
      RECT  55.0 12.55 55.29 12.84 ;
      RECT  54.65 12.53 54.79 13.06 ;
      RECT  53.55 12.04 53.84 12.26 ;
      RECT  52.83 11.9 53.11 12.0 ;
      RECT  52.69 9.47 55.77 9.64 ;
      RECT  53.69 12.33 53.86 12.35 ;
      RECT  52.84 10.44 53.15 10.73 ;
      RECT  49.61 11.73 52.69 11.9 ;
      RECT  52.69 11.73 55.77 11.9 ;
      RECT  42.55 9.485 55.77 9.625 ;
      RECT  50.96 2.08 51.61 2.23 ;
      RECT  49.98 0.09 50.15 0.52 ;
      RECT  50.81 4.93 51.1 5.22 ;
      RECT  51.48 0.56 51.81 1.07 ;
      RECT  51.87 2.59 52.2 2.67 ;
      RECT  50.3 6.93 50.59 6.99 ;
      RECT  51.34 1.47 51.63 1.76 ;
      RECT  51.87 2.84 52.2 2.92 ;
      RECT  50.49 1.45 50.97 1.8 ;
      RECT  49.81 2.23 50.1 2.29 ;
      RECT  49.61 5.66 52.69 5.83 ;
      RECT  50.86 3.56 51.01 4.2 ;
      RECT  49.92 0.52 50.21 1.24 ;
      RECT  49.61 -0.08 52.69 0.09 ;
      RECT  50.81 2.46 51.1 2.52 ;
      RECT  51.44 -0.17 51.79 -0.08 ;
      RECT  50.81 3.27 51.1 3.56 ;
      RECT  49.79 6.14 50.12 6.22 ;
      RECT  51.52 4.37 51.87 4.46 ;
      RECT  50.86 4.37 51.01 4.93 ;
      RECT  51.48 1.07 52.48 1.27 ;
      RECT  50.64 0.53 50.97 1.45 ;
      RECT  49.61 2.67 52.69 2.84 ;
      RECT  52.19 0.09 52.36 0.5 ;
      RECT  50.81 6.39 51.1 6.45 ;
      RECT  50.81 6.16 51.1 6.22 ;
      RECT  50.81 2.23 51.1 2.29 ;
      RECT  49.76 1.45 50.11 1.8 ;
      RECT  51.46 1.76 51.61 2.08 ;
      RECT  52.13 1.27 52.48 1.31 ;
      RECT  49.77 6.48 50.12 6.83 ;
      RECT  50.3 7.15 52.69 7.16 ;
      RECT  49.97 5.6 50.26 5.66 ;
      RECT  52.13 0.5 52.42 0.79 ;
      RECT  51.36 7.16 51.71 7.25 ;
      RECT  51.44 0.09 51.79 0.18 ;
      RECT  49.61 6.99 52.69 7.15 ;
      RECT  51.52 4.11 51.87 4.2 ;
      RECT  52.13 0.96 52.48 1.07 ;
      RECT  50.3 7.16 50.59 7.22 ;
      RECT  51.36 6.9 51.71 6.99 ;
      RECT  49.79 6.39 50.12 6.48 ;
      RECT  49.61 4.2 52.69 4.37 ;
      RECT  49.81 2.29 51.1 2.46 ;
      RECT  49.81 2.46 50.1 2.52 ;
      RECT  49.79 6.22 51.1 6.39 ;
      RECT  52.11 6.46 52.28 6.99 ;
      RECT  49.97 5.83 50.26 5.89 ;
      RECT  52.05 6.17 52.34 6.46 ;
      RECT  54.04 2.08 54.69 2.23 ;
      RECT  53.06 0.09 53.23 0.52 ;
      RECT  53.89 4.93 54.18 5.22 ;
      RECT  54.56 0.56 54.89 1.07 ;
      RECT  54.95 2.59 55.28 2.67 ;
      RECT  53.38 6.93 53.67 6.99 ;
      RECT  54.42 1.47 54.71 1.76 ;
      RECT  54.95 2.84 55.28 2.92 ;
      RECT  53.57 1.45 54.05 1.8 ;
      RECT  52.89 2.23 53.18 2.29 ;
      RECT  52.69 5.66 55.77 5.83 ;
      RECT  53.94 3.56 54.09 4.2 ;
      RECT  53.0 0.52 53.29 1.24 ;
      RECT  52.69 -0.08 55.77 0.09 ;
      RECT  53.89 2.46 54.18 2.52 ;
      RECT  54.52 -0.17 54.87 -0.08 ;
      RECT  53.89 3.27 54.18 3.56 ;
      RECT  52.87 6.14 53.2 6.22 ;
      RECT  54.6 4.37 54.95 4.46 ;
      RECT  53.94 4.37 54.09 4.93 ;
      RECT  54.56 1.07 55.56 1.27 ;
      RECT  53.72 0.53 54.05 1.45 ;
      RECT  52.69 2.67 55.77 2.84 ;
      RECT  55.27 0.09 55.44 0.5 ;
      RECT  53.89 6.39 54.18 6.45 ;
      RECT  53.89 6.16 54.18 6.22 ;
      RECT  53.89 2.23 54.18 2.29 ;
      RECT  52.84 1.45 53.19 1.8 ;
      RECT  54.54 1.76 54.69 2.08 ;
      RECT  55.21 1.27 55.56 1.31 ;
      RECT  52.85 6.48 53.2 6.83 ;
      RECT  53.38 7.15 55.77 7.16 ;
      RECT  53.05 5.6 53.34 5.66 ;
      RECT  55.21 0.5 55.5 0.79 ;
      RECT  54.44 7.16 54.79 7.25 ;
      RECT  54.52 0.09 54.87 0.18 ;
      RECT  52.69 6.99 55.77 7.15 ;
      RECT  54.6 4.11 54.95 4.2 ;
      RECT  55.21 0.96 55.56 1.07 ;
      RECT  53.38 7.16 53.67 7.22 ;
      RECT  54.44 6.9 54.79 6.99 ;
      RECT  52.87 6.39 53.2 6.48 ;
      RECT  52.69 4.2 55.77 4.37 ;
      RECT  52.89 2.29 54.18 2.46 ;
      RECT  52.89 2.46 53.18 2.52 ;
      RECT  52.87 6.22 54.18 6.39 ;
      RECT  55.19 6.46 55.36 6.99 ;
      RECT  53.05 5.83 53.34 5.89 ;
      RECT  55.13 6.17 55.42 6.46 ;
      RECT  49.61 2.67 52.69 2.84 ;
      RECT  52.69 2.67 55.77 2.84 ;
      RECT  42.55 5.66 55.77 5.8 ;
      RECT  49.61 11.9 52.69 11.73 ;
      RECT  52.69 11.9 55.77 11.73 ;
      RECT  49.61 2.84 52.69 2.67 ;
      RECT  52.69 2.84 55.77 2.67 ;
      RECT  42.55 9.625 55.77 9.485 ;
      RECT  42.55 16.925 55.77 16.785 ;
      RECT  42.55 5.8 55.77 5.66 ;
      RECT  49.61 11.73 52.69 11.9 ;
      RECT  52.69 11.73 55.77 11.9 ;
      RECT  49.61 2.67 52.69 2.84 ;
      RECT  52.69 2.67 55.77 2.84 ;
      RECT  -52.26 -7.44 -47.34 -7.19 ;
      RECT  -55.37 -7.8 -54.69 -7.48 ;
      RECT  -46.46 -6.74 -46.13 -6.62 ;
      RECT  -54.5 -7.92 -54.21 -7.89 ;
      RECT  -55.45 -9.48 -42.92 -9.15 ;
      RECT  -47.54 -7.61 -47.34 -7.44 ;
      RECT  -54.5 -7.69 -54.21 -7.63 ;
      RECT  -46.85 -7.84 -46.55 -7.73 ;
      RECT  -47.54 -6.94 -46.13 -6.74 ;
      RECT  -52.26 -6.95 -51.93 -6.94 ;
      RECT  -48.18 -6.95 -47.85 -6.94 ;
      RECT  -54.22 -6.98 -53.59 -6.66 ;
      RECT  -47.58 -7.94 -47.25 -7.61 ;
      RECT  -53.34 -6.94 -47.85 -6.74 ;
      RECT  -52.65 -8.05 -49.36 -7.84 ;
      RECT  -49.69 -8.1 -49.36 -8.05 ;
      RECT  -48.18 -6.74 -47.85 -6.62 ;
      RECT  -52.26 -6.74 -51.93 -6.62 ;
      RECT  -53.38 -7.69 -53.05 -7.61 ;
      RECT  -52.65 -7.84 -52.35 -7.74 ;
      RECT  -43.66 -7.84 -43.32 -7.81 ;
      RECT  -46.85 -8.04 -43.32 -7.84 ;
      RECT  -49.69 -7.84 -49.36 -7.77 ;
      RECT  -45.32 -7.29 -44.69 -6.97 ;
      RECT  -52.26 -7.19 -51.93 -7.16 ;
      RECT  -53.38 -7.94 -53.05 -7.89 ;
      RECT  -43.66 -8.14 -43.32 -8.04 ;
      RECT  -46.46 -6.95 -46.13 -6.94 ;
      RECT  -52.26 -7.49 -51.93 -7.44 ;
      RECT  -54.5 -7.89 -53.05 -7.69 ;
      RECT  -55.39 -5.39 -42.74 -5.06 ;
      RECT  -53.34 -7.61 -53.14 -6.94 ;
      RECT  -47.54 -7.19 -47.34 -6.94 ;
      RECT  -55.39 -5.39 -31.52 -5.06 ;
      RECT  -55.45 -9.48 -31.58 -9.15 ;
      RECT  -52.26 -3.0 -47.34 -3.25 ;
      RECT  -55.37 -2.64 -54.69 -2.96 ;
      RECT  -46.46 -3.7 -46.13 -3.82 ;
      RECT  -54.5 -2.52 -54.21 -2.55 ;
      RECT  -55.45 -0.96 -42.92 -1.29 ;
      RECT  -47.54 -2.83 -47.34 -3.0 ;
      RECT  -54.5 -2.75 -54.21 -2.81 ;
      RECT  -46.85 -2.6 -46.55 -2.71 ;
      RECT  -47.54 -3.5 -46.13 -3.7 ;
      RECT  -52.26 -3.49 -51.93 -3.5 ;
      RECT  -48.18 -3.49 -47.85 -3.5 ;
      RECT  -54.22 -3.46 -53.59 -3.78 ;
      RECT  -47.58 -2.5 -47.25 -2.83 ;
      RECT  -53.34 -3.5 -47.85 -3.7 ;
      RECT  -52.65 -2.39 -49.36 -2.6 ;
      RECT  -49.69 -2.34 -49.36 -2.39 ;
      RECT  -48.18 -3.7 -47.85 -3.82 ;
      RECT  -52.26 -3.7 -51.93 -3.82 ;
      RECT  -53.38 -2.75 -53.05 -2.83 ;
      RECT  -52.65 -2.6 -52.35 -2.7 ;
      RECT  -43.66 -2.6 -43.32 -2.63 ;
      RECT  -46.85 -2.4 -43.32 -2.6 ;
      RECT  -49.69 -2.6 -49.36 -2.67 ;
      RECT  -45.32 -3.15 -44.69 -3.47 ;
      RECT  -52.26 -3.25 -51.93 -3.28 ;
      RECT  -53.38 -2.5 -53.05 -2.55 ;
      RECT  -43.66 -2.3 -43.32 -2.4 ;
      RECT  -46.46 -3.49 -46.13 -3.5 ;
      RECT  -52.26 -2.95 -51.93 -3.0 ;
      RECT  -54.5 -2.55 -53.05 -2.75 ;
      RECT  -55.39 -5.05 -42.74 -5.38 ;
      RECT  -53.34 -2.83 -53.14 -3.5 ;
      RECT  -47.54 -3.25 -47.34 -3.5 ;
      RECT  -55.39 -5.05 -31.52 -5.38 ;
      RECT  -55.45 -0.96 -31.58 -1.29 ;
      RECT  -10.84 103.28 -5.92 103.53 ;
      RECT  -13.95 102.92 -13.27 103.24 ;
      RECT  -5.04 103.98 -4.71 104.1 ;
      RECT  -13.08 102.8 -12.79 102.83 ;
      RECT  -14.03 101.24 -1.5 101.57 ;
      RECT  -6.12 103.11 -5.92 103.28 ;
      RECT  -13.08 103.03 -12.79 103.09 ;
      RECT  -5.43 102.88 -5.13 102.99 ;
      RECT  -6.12 103.78 -4.71 103.98 ;
      RECT  -10.84 103.77 -10.51 103.78 ;
      RECT  -6.76 103.77 -6.43 103.78 ;
      RECT  -12.8 103.74 -12.17 104.06 ;
      RECT  -6.16 102.78 -5.83 103.11 ;
      RECT  -11.92 103.78 -6.43 103.98 ;
      RECT  -11.23 102.67 -7.94 102.88 ;
      RECT  -8.27 102.62 -7.94 102.67 ;
      RECT  -6.76 103.98 -6.43 104.1 ;
      RECT  -10.84 103.98 -10.51 104.1 ;
      RECT  -11.96 103.03 -11.63 103.11 ;
      RECT  -11.23 102.88 -10.93 102.98 ;
      RECT  -2.24 102.88 -1.9 102.91 ;
      RECT  -5.43 102.68 -1.9 102.88 ;
      RECT  -8.27 102.88 -7.94 102.95 ;
      RECT  -3.9 103.43 -3.27 103.75 ;
      RECT  -10.84 103.53 -10.51 103.56 ;
      RECT  -11.96 102.78 -11.63 102.83 ;
      RECT  -2.24 102.58 -1.9 102.68 ;
      RECT  -5.04 103.77 -4.71 103.78 ;
      RECT  -10.84 103.23 -10.51 103.28 ;
      RECT  -13.08 102.83 -11.63 103.03 ;
      RECT  -13.97 105.33 -1.32 105.66 ;
      RECT  -11.92 103.11 -11.72 103.78 ;
      RECT  -6.12 103.53 -5.92 103.78 ;
      RECT  -10.84 107.72 -5.92 107.47 ;
      RECT  -13.95 108.08 -13.27 107.76 ;
      RECT  -5.04 107.02 -4.71 106.9 ;
      RECT  -13.08 108.2 -12.79 108.17 ;
      RECT  -14.03 109.76 -1.5 109.43 ;
      RECT  -6.12 107.89 -5.92 107.72 ;
      RECT  -13.08 107.97 -12.79 107.91 ;
      RECT  -5.43 108.12 -5.13 108.01 ;
      RECT  -6.12 107.22 -4.71 107.02 ;
      RECT  -10.84 107.23 -10.51 107.22 ;
      RECT  -6.76 107.23 -6.43 107.22 ;
      RECT  -12.8 107.26 -12.17 106.94 ;
      RECT  -6.16 108.22 -5.83 107.89 ;
      RECT  -11.92 107.22 -6.43 107.02 ;
      RECT  -11.23 108.33 -7.94 108.12 ;
      RECT  -8.27 108.38 -7.94 108.33 ;
      RECT  -6.76 107.02 -6.43 106.9 ;
      RECT  -10.84 107.02 -10.51 106.9 ;
      RECT  -11.96 107.97 -11.63 107.89 ;
      RECT  -11.23 108.12 -10.93 108.02 ;
      RECT  -2.24 108.12 -1.9 108.09 ;
      RECT  -5.43 108.32 -1.9 108.12 ;
      RECT  -8.27 108.12 -7.94 108.05 ;
      RECT  -3.9 107.57 -3.27 107.25 ;
      RECT  -10.84 107.47 -10.51 107.44 ;
      RECT  -11.96 108.22 -11.63 108.17 ;
      RECT  -2.24 108.42 -1.9 108.32 ;
      RECT  -5.04 107.23 -4.71 107.22 ;
      RECT  -10.84 107.77 -10.51 107.72 ;
      RECT  -13.08 108.17 -11.63 107.97 ;
      RECT  -13.97 105.67 -1.32 105.34 ;
      RECT  -11.92 107.89 -11.72 107.22 ;
      RECT  -6.12 107.47 -5.92 107.22 ;
      RECT  -10.84 111.46 -5.92 111.71 ;
      RECT  -13.95 111.1 -13.27 111.42 ;
      RECT  -5.04 112.16 -4.71 112.28 ;
      RECT  -13.08 110.98 -12.79 111.01 ;
      RECT  -14.03 109.42 -1.5 109.75 ;
      RECT  -6.12 111.29 -5.92 111.46 ;
      RECT  -13.08 111.21 -12.79 111.27 ;
      RECT  -5.43 111.06 -5.13 111.17 ;
      RECT  -6.12 111.96 -4.71 112.16 ;
      RECT  -10.84 111.95 -10.51 111.96 ;
      RECT  -6.76 111.95 -6.43 111.96 ;
      RECT  -12.8 111.92 -12.17 112.24 ;
      RECT  -6.16 110.96 -5.83 111.29 ;
      RECT  -11.92 111.96 -6.43 112.16 ;
      RECT  -11.23 110.85 -7.94 111.06 ;
      RECT  -8.27 110.8 -7.94 110.85 ;
      RECT  -6.76 112.16 -6.43 112.28 ;
      RECT  -10.84 112.16 -10.51 112.28 ;
      RECT  -11.96 111.21 -11.63 111.29 ;
      RECT  -11.23 111.06 -10.93 111.16 ;
      RECT  -2.24 111.06 -1.9 111.09 ;
      RECT  -5.43 110.86 -1.9 111.06 ;
      RECT  -8.27 111.06 -7.94 111.13 ;
      RECT  -3.9 111.61 -3.27 111.93 ;
      RECT  -10.84 111.71 -10.51 111.74 ;
      RECT  -11.96 110.96 -11.63 111.01 ;
      RECT  -2.24 110.76 -1.9 110.86 ;
      RECT  -5.04 111.95 -4.71 111.96 ;
      RECT  -10.84 111.41 -10.51 111.46 ;
      RECT  -13.08 111.01 -11.63 111.21 ;
      RECT  -13.97 113.51 -1.32 113.84 ;
      RECT  -11.92 111.29 -11.72 111.96 ;
      RECT  -6.12 111.71 -5.92 111.96 ;
      RECT  -10.84 115.9 -5.92 115.65 ;
      RECT  -13.95 116.26 -13.27 115.94 ;
      RECT  -5.04 115.2 -4.71 115.08 ;
      RECT  -13.08 116.38 -12.79 116.35 ;
      RECT  -14.03 117.94 -1.5 117.61 ;
      RECT  -6.12 116.07 -5.92 115.9 ;
      RECT  -13.08 116.15 -12.79 116.09 ;
      RECT  -5.43 116.3 -5.13 116.19 ;
      RECT  -6.12 115.4 -4.71 115.2 ;
      RECT  -10.84 115.41 -10.51 115.4 ;
      RECT  -6.76 115.41 -6.43 115.4 ;
      RECT  -12.8 115.44 -12.17 115.12 ;
      RECT  -6.16 116.4 -5.83 116.07 ;
      RECT  -11.92 115.4 -6.43 115.2 ;
      RECT  -11.23 116.51 -7.94 116.3 ;
      RECT  -8.27 116.56 -7.94 116.51 ;
      RECT  -6.76 115.2 -6.43 115.08 ;
      RECT  -10.84 115.2 -10.51 115.08 ;
      RECT  -11.96 116.15 -11.63 116.07 ;
      RECT  -11.23 116.3 -10.93 116.2 ;
      RECT  -2.24 116.3 -1.9 116.27 ;
      RECT  -5.43 116.5 -1.9 116.3 ;
      RECT  -8.27 116.3 -7.94 116.23 ;
      RECT  -3.9 115.75 -3.27 115.43 ;
      RECT  -10.84 115.65 -10.51 115.62 ;
      RECT  -11.96 116.4 -11.63 116.35 ;
      RECT  -2.24 116.6 -1.9 116.5 ;
      RECT  -5.04 115.41 -4.71 115.4 ;
      RECT  -10.84 115.95 -10.51 115.9 ;
      RECT  -13.08 116.35 -11.63 116.15 ;
      RECT  -13.97 113.85 -1.32 113.52 ;
      RECT  -11.92 116.07 -11.72 115.4 ;
      RECT  -6.12 115.65 -5.92 115.4 ;
      RECT  14.58 -7.44 19.5 -7.19 ;
      RECT  11.47 -7.8 12.15 -7.48 ;
      RECT  20.38 -6.74 20.71 -6.62 ;
      RECT  12.34 -7.92 12.63 -7.89 ;
      RECT  11.39 -9.48 23.92 -9.15 ;
      RECT  19.3 -7.61 19.5 -7.44 ;
      RECT  12.34 -7.69 12.63 -7.63 ;
      RECT  19.99 -7.84 20.29 -7.73 ;
      RECT  19.3 -6.94 20.71 -6.74 ;
      RECT  14.58 -6.95 14.91 -6.94 ;
      RECT  18.66 -6.95 18.99 -6.94 ;
      RECT  12.62 -6.98 13.25 -6.66 ;
      RECT  19.26 -7.94 19.59 -7.61 ;
      RECT  13.5 -6.94 18.99 -6.74 ;
      RECT  14.19 -8.05 17.48 -7.84 ;
      RECT  17.15 -8.1 17.48 -8.05 ;
      RECT  18.66 -6.74 18.99 -6.62 ;
      RECT  14.58 -6.74 14.91 -6.62 ;
      RECT  13.46 -7.69 13.79 -7.61 ;
      RECT  14.19 -7.84 14.49 -7.74 ;
      RECT  23.18 -7.84 23.52 -7.81 ;
      RECT  19.99 -8.04 23.52 -7.84 ;
      RECT  17.15 -7.84 17.48 -7.77 ;
      RECT  21.52 -7.29 22.15 -6.97 ;
      RECT  14.58 -7.19 14.91 -7.16 ;
      RECT  13.46 -7.94 13.79 -7.89 ;
      RECT  23.18 -8.14 23.52 -8.04 ;
      RECT  20.38 -6.95 20.71 -6.94 ;
      RECT  14.58 -7.49 14.91 -7.44 ;
      RECT  12.34 -7.89 13.79 -7.69 ;
      RECT  11.45 -5.39 24.1 -5.06 ;
      RECT  13.5 -7.61 13.7 -6.94 ;
      RECT  19.3 -7.19 19.5 -6.94 ;
      RECT  27.29 -7.44 32.21 -7.19 ;
      RECT  24.18 -7.8 24.86 -7.48 ;
      RECT  33.09 -6.74 33.42 -6.62 ;
      RECT  25.05 -7.92 25.34 -7.89 ;
      RECT  24.1 -9.48 36.63 -9.15 ;
      RECT  32.01 -7.61 32.21 -7.44 ;
      RECT  25.05 -7.69 25.34 -7.63 ;
      RECT  32.7 -7.84 33.0 -7.73 ;
      RECT  32.01 -6.94 33.42 -6.74 ;
      RECT  27.29 -6.95 27.62 -6.94 ;
      RECT  31.37 -6.95 31.7 -6.94 ;
      RECT  25.33 -6.98 25.96 -6.66 ;
      RECT  31.97 -7.94 32.3 -7.61 ;
      RECT  26.21 -6.94 31.7 -6.74 ;
      RECT  26.9 -8.05 30.19 -7.84 ;
      RECT  29.86 -8.1 30.19 -8.05 ;
      RECT  31.37 -6.74 31.7 -6.62 ;
      RECT  27.29 -6.74 27.62 -6.62 ;
      RECT  26.17 -7.69 26.5 -7.61 ;
      RECT  26.9 -7.84 27.2 -7.74 ;
      RECT  35.89 -7.84 36.23 -7.81 ;
      RECT  32.7 -8.04 36.23 -7.84 ;
      RECT  29.86 -7.84 30.19 -7.77 ;
      RECT  34.23 -7.29 34.86 -6.97 ;
      RECT  27.29 -7.19 27.62 -7.16 ;
      RECT  26.17 -7.94 26.5 -7.89 ;
      RECT  35.89 -8.14 36.23 -8.04 ;
      RECT  33.09 -6.95 33.42 -6.94 ;
      RECT  27.29 -7.49 27.62 -7.44 ;
      RECT  25.05 -7.89 26.5 -7.69 ;
      RECT  24.16 -5.39 36.81 -5.06 ;
      RECT  26.21 -7.61 26.41 -6.94 ;
      RECT  32.01 -7.19 32.21 -6.94 ;
   LAYER  m2 ;
      RECT  50.97 33.07 51.11 34.06 ;
      RECT  51.85 35.73 51.99 37.99 ;
      RECT  50.97 34.06 51.32 34.41 ;
      RECT  50.01 33.09 50.46 33.54 ;
      RECT  50.01 37.32 50.46 37.77 ;
      RECT  51.85 33.07 51.99 35.38 ;
      RECT  50.97 34.41 51.11 37.99 ;
      RECT  51.76 35.38 52.11 35.73 ;
      RECT  50.97 42.25 51.11 41.26 ;
      RECT  51.85 39.59 51.99 37.33 ;
      RECT  50.97 41.26 51.32 40.91 ;
      RECT  50.01 42.23 50.46 41.78 ;
      RECT  50.01 38.0 50.46 37.55 ;
      RECT  51.85 42.25 51.99 39.94 ;
      RECT  50.97 40.91 51.11 37.33 ;
      RECT  51.76 39.94 52.11 39.59 ;
      RECT  50.97 41.77 51.11 42.76 ;
      RECT  51.85 44.43 51.99 46.69 ;
      RECT  50.97 42.76 51.32 43.11 ;
      RECT  50.01 41.79 50.46 42.24 ;
      RECT  50.01 46.02 50.46 46.47 ;
      RECT  51.85 41.77 51.99 44.08 ;
      RECT  50.97 43.11 51.11 46.69 ;
      RECT  51.76 44.08 52.11 44.43 ;
      RECT  50.97 50.95 51.11 49.96 ;
      RECT  51.85 48.29 51.99 46.03 ;
      RECT  50.97 49.96 51.32 49.61 ;
      RECT  50.01 50.93 50.46 50.48 ;
      RECT  50.01 46.7 50.46 46.25 ;
      RECT  51.85 50.95 51.99 48.64 ;
      RECT  50.97 49.61 51.11 46.03 ;
      RECT  51.76 48.64 52.11 48.29 ;
      RECT  50.97 50.47 51.11 51.46 ;
      RECT  51.85 53.13 51.99 55.39 ;
      RECT  50.97 51.46 51.32 51.81 ;
      RECT  50.01 50.49 50.46 50.94 ;
      RECT  50.01 54.72 50.46 55.17 ;
      RECT  51.85 50.47 51.99 52.78 ;
      RECT  50.97 51.81 51.11 55.39 ;
      RECT  51.76 52.78 52.11 53.13 ;
      RECT  50.97 59.65 51.11 58.66 ;
      RECT  51.85 56.99 51.99 54.73 ;
      RECT  50.97 58.66 51.32 58.31 ;
      RECT  50.01 59.63 50.46 59.18 ;
      RECT  50.01 55.4 50.46 54.95 ;
      RECT  51.85 59.65 51.99 57.34 ;
      RECT  50.97 58.31 51.11 54.73 ;
      RECT  51.76 57.34 52.11 56.99 ;
      RECT  50.97 59.17 51.11 60.16 ;
      RECT  51.85 61.83 51.99 64.09 ;
      RECT  50.97 60.16 51.32 60.51 ;
      RECT  50.01 59.19 50.46 59.64 ;
      RECT  50.01 63.42 50.46 63.87 ;
      RECT  51.85 59.17 51.99 61.48 ;
      RECT  50.97 60.51 51.11 64.09 ;
      RECT  51.76 61.48 52.11 61.83 ;
      RECT  50.97 68.35 51.11 67.36 ;
      RECT  51.85 65.69 51.99 63.43 ;
      RECT  50.97 67.36 51.32 67.01 ;
      RECT  50.01 68.33 50.46 67.88 ;
      RECT  50.01 64.1 50.46 63.65 ;
      RECT  51.85 68.35 51.99 66.04 ;
      RECT  50.97 67.01 51.11 63.43 ;
      RECT  51.76 66.04 52.11 65.69 ;
      RECT  50.97 67.87 51.11 68.86 ;
      RECT  51.85 70.53 51.99 72.79 ;
      RECT  50.97 68.86 51.32 69.21 ;
      RECT  50.01 67.89 50.46 68.34 ;
      RECT  50.01 72.12 50.46 72.57 ;
      RECT  51.85 67.87 51.99 70.18 ;
      RECT  50.97 69.21 51.11 72.79 ;
      RECT  51.76 70.18 52.11 70.53 ;
      RECT  50.97 77.05 51.11 76.06 ;
      RECT  51.85 74.39 51.99 72.13 ;
      RECT  50.97 76.06 51.32 75.71 ;
      RECT  50.01 77.03 50.46 76.58 ;
      RECT  50.01 72.8 50.46 72.35 ;
      RECT  51.85 77.05 51.99 74.74 ;
      RECT  50.97 75.71 51.11 72.13 ;
      RECT  51.76 74.74 52.11 74.39 ;
      RECT  50.97 76.57 51.11 77.56 ;
      RECT  51.85 79.23 51.99 81.49 ;
      RECT  50.97 77.56 51.32 77.91 ;
      RECT  50.01 76.59 50.46 77.04 ;
      RECT  50.01 80.82 50.46 81.27 ;
      RECT  51.85 76.57 51.99 78.88 ;
      RECT  50.97 77.91 51.11 81.49 ;
      RECT  51.76 78.88 52.11 79.23 ;
      RECT  50.97 85.75 51.11 84.76 ;
      RECT  51.85 83.09 51.99 80.83 ;
      RECT  50.97 84.76 51.32 84.41 ;
      RECT  50.01 85.73 50.46 85.28 ;
      RECT  50.01 81.5 50.46 81.05 ;
      RECT  51.85 85.75 51.99 83.44 ;
      RECT  50.97 84.41 51.11 80.83 ;
      RECT  51.76 83.44 52.11 83.09 ;
      RECT  50.97 85.27 51.11 86.26 ;
      RECT  51.85 87.93 51.99 90.19 ;
      RECT  50.97 86.26 51.32 86.61 ;
      RECT  50.01 85.29 50.46 85.74 ;
      RECT  50.01 89.52 50.46 89.97 ;
      RECT  51.85 85.27 51.99 87.58 ;
      RECT  50.97 86.61 51.11 90.19 ;
      RECT  51.76 87.58 52.11 87.93 ;
      RECT  50.97 94.45 51.11 93.46 ;
      RECT  51.85 91.79 51.99 89.53 ;
      RECT  50.97 93.46 51.32 93.11 ;
      RECT  50.01 94.43 50.46 93.98 ;
      RECT  50.01 90.2 50.46 89.75 ;
      RECT  51.85 94.45 51.99 92.14 ;
      RECT  50.97 93.11 51.11 89.53 ;
      RECT  51.76 92.14 52.11 91.79 ;
      RECT  50.97 93.97 51.11 94.96 ;
      RECT  51.85 96.63 51.99 98.89 ;
      RECT  50.97 94.96 51.32 95.31 ;
      RECT  50.01 93.99 50.46 94.44 ;
      RECT  50.01 98.22 50.46 98.67 ;
      RECT  51.85 93.97 51.99 96.28 ;
      RECT  50.97 95.31 51.11 98.89 ;
      RECT  51.76 96.28 52.11 96.63 ;
      RECT  50.97 103.15 51.11 102.16 ;
      RECT  51.85 100.49 51.99 98.23 ;
      RECT  50.97 102.16 51.32 101.81 ;
      RECT  50.01 103.13 50.46 102.68 ;
      RECT  50.01 98.9 50.46 98.45 ;
      RECT  51.85 103.15 51.99 100.84 ;
      RECT  50.97 101.81 51.11 98.23 ;
      RECT  51.76 100.84 52.11 100.49 ;
      RECT  54.05 33.07 54.19 34.06 ;
      RECT  54.93 35.73 55.07 37.99 ;
      RECT  54.05 34.06 54.4 34.41 ;
      RECT  53.09 33.09 53.54 33.54 ;
      RECT  53.09 37.32 53.54 37.77 ;
      RECT  54.93 33.07 55.07 35.38 ;
      RECT  54.05 34.41 54.19 37.99 ;
      RECT  54.84 35.38 55.19 35.73 ;
      RECT  54.05 42.25 54.19 41.26 ;
      RECT  54.93 39.59 55.07 37.33 ;
      RECT  54.05 41.26 54.4 40.91 ;
      RECT  53.09 42.23 53.54 41.78 ;
      RECT  53.09 38.0 53.54 37.55 ;
      RECT  54.93 42.25 55.07 39.94 ;
      RECT  54.05 40.91 54.19 37.33 ;
      RECT  54.84 39.94 55.19 39.59 ;
      RECT  54.05 41.77 54.19 42.76 ;
      RECT  54.93 44.43 55.07 46.69 ;
      RECT  54.05 42.76 54.4 43.11 ;
      RECT  53.09 41.79 53.54 42.24 ;
      RECT  53.09 46.02 53.54 46.47 ;
      RECT  54.93 41.77 55.07 44.08 ;
      RECT  54.05 43.11 54.19 46.69 ;
      RECT  54.84 44.08 55.19 44.43 ;
      RECT  54.05 50.95 54.19 49.96 ;
      RECT  54.93 48.29 55.07 46.03 ;
      RECT  54.05 49.96 54.4 49.61 ;
      RECT  53.09 50.93 53.54 50.48 ;
      RECT  53.09 46.7 53.54 46.25 ;
      RECT  54.93 50.95 55.07 48.64 ;
      RECT  54.05 49.61 54.19 46.03 ;
      RECT  54.84 48.64 55.19 48.29 ;
      RECT  54.05 50.47 54.19 51.46 ;
      RECT  54.93 53.13 55.07 55.39 ;
      RECT  54.05 51.46 54.4 51.81 ;
      RECT  53.09 50.49 53.54 50.94 ;
      RECT  53.09 54.72 53.54 55.17 ;
      RECT  54.93 50.47 55.07 52.78 ;
      RECT  54.05 51.81 54.19 55.39 ;
      RECT  54.84 52.78 55.19 53.13 ;
      RECT  54.05 59.65 54.19 58.66 ;
      RECT  54.93 56.99 55.07 54.73 ;
      RECT  54.05 58.66 54.4 58.31 ;
      RECT  53.09 59.63 53.54 59.18 ;
      RECT  53.09 55.4 53.54 54.95 ;
      RECT  54.93 59.65 55.07 57.34 ;
      RECT  54.05 58.31 54.19 54.73 ;
      RECT  54.84 57.34 55.19 56.99 ;
      RECT  54.05 59.17 54.19 60.16 ;
      RECT  54.93 61.83 55.07 64.09 ;
      RECT  54.05 60.16 54.4 60.51 ;
      RECT  53.09 59.19 53.54 59.64 ;
      RECT  53.09 63.42 53.54 63.87 ;
      RECT  54.93 59.17 55.07 61.48 ;
      RECT  54.05 60.51 54.19 64.09 ;
      RECT  54.84 61.48 55.19 61.83 ;
      RECT  54.05 68.35 54.19 67.36 ;
      RECT  54.93 65.69 55.07 63.43 ;
      RECT  54.05 67.36 54.4 67.01 ;
      RECT  53.09 68.33 53.54 67.88 ;
      RECT  53.09 64.1 53.54 63.65 ;
      RECT  54.93 68.35 55.07 66.04 ;
      RECT  54.05 67.01 54.19 63.43 ;
      RECT  54.84 66.04 55.19 65.69 ;
      RECT  54.05 67.87 54.19 68.86 ;
      RECT  54.93 70.53 55.07 72.79 ;
      RECT  54.05 68.86 54.4 69.21 ;
      RECT  53.09 67.89 53.54 68.34 ;
      RECT  53.09 72.12 53.54 72.57 ;
      RECT  54.93 67.87 55.07 70.18 ;
      RECT  54.05 69.21 54.19 72.79 ;
      RECT  54.84 70.18 55.19 70.53 ;
      RECT  54.05 77.05 54.19 76.06 ;
      RECT  54.93 74.39 55.07 72.13 ;
      RECT  54.05 76.06 54.4 75.71 ;
      RECT  53.09 77.03 53.54 76.58 ;
      RECT  53.09 72.8 53.54 72.35 ;
      RECT  54.93 77.05 55.07 74.74 ;
      RECT  54.05 75.71 54.19 72.13 ;
      RECT  54.84 74.74 55.19 74.39 ;
      RECT  54.05 76.57 54.19 77.56 ;
      RECT  54.93 79.23 55.07 81.49 ;
      RECT  54.05 77.56 54.4 77.91 ;
      RECT  53.09 76.59 53.54 77.04 ;
      RECT  53.09 80.82 53.54 81.27 ;
      RECT  54.93 76.57 55.07 78.88 ;
      RECT  54.05 77.91 54.19 81.49 ;
      RECT  54.84 78.88 55.19 79.23 ;
      RECT  54.05 85.75 54.19 84.76 ;
      RECT  54.93 83.09 55.07 80.83 ;
      RECT  54.05 84.76 54.4 84.41 ;
      RECT  53.09 85.73 53.54 85.28 ;
      RECT  53.09 81.5 53.54 81.05 ;
      RECT  54.93 85.75 55.07 83.44 ;
      RECT  54.05 84.41 54.19 80.83 ;
      RECT  54.84 83.44 55.19 83.09 ;
      RECT  54.05 85.27 54.19 86.26 ;
      RECT  54.93 87.93 55.07 90.19 ;
      RECT  54.05 86.26 54.4 86.61 ;
      RECT  53.09 85.29 53.54 85.74 ;
      RECT  53.09 89.52 53.54 89.97 ;
      RECT  54.93 85.27 55.07 87.58 ;
      RECT  54.05 86.61 54.19 90.19 ;
      RECT  54.84 87.58 55.19 87.93 ;
      RECT  54.05 94.45 54.19 93.46 ;
      RECT  54.93 91.79 55.07 89.53 ;
      RECT  54.05 93.46 54.4 93.11 ;
      RECT  53.09 94.43 53.54 93.98 ;
      RECT  53.09 90.2 53.54 89.75 ;
      RECT  54.93 94.45 55.07 92.14 ;
      RECT  54.05 93.11 54.19 89.53 ;
      RECT  54.84 92.14 55.19 91.79 ;
      RECT  54.05 93.97 54.19 94.96 ;
      RECT  54.93 96.63 55.07 98.89 ;
      RECT  54.05 94.96 54.4 95.31 ;
      RECT  53.09 93.99 53.54 94.44 ;
      RECT  53.09 98.22 53.54 98.67 ;
      RECT  54.93 93.97 55.07 96.28 ;
      RECT  54.05 95.31 54.19 98.89 ;
      RECT  54.84 96.28 55.19 96.63 ;
      RECT  54.05 103.15 54.19 102.16 ;
      RECT  54.93 100.49 55.07 98.23 ;
      RECT  54.05 102.16 54.4 101.81 ;
      RECT  53.09 103.13 53.54 102.68 ;
      RECT  53.09 98.9 53.54 98.45 ;
      RECT  54.93 103.15 55.07 100.84 ;
      RECT  54.05 101.81 54.19 98.23 ;
      RECT  54.84 100.84 55.19 100.49 ;
      RECT  50.97 33.31 51.32 102.91 ;
      RECT  51.76 33.31 52.11 102.91 ;
      RECT  54.05 33.31 54.4 102.91 ;
      RECT  54.84 33.31 55.19 102.91 ;
      RECT  47.89 24.37 48.03 25.36 ;
      RECT  48.77 27.03 48.91 29.29 ;
      RECT  47.89 25.36 48.24 25.71 ;
      RECT  46.93 24.39 47.38 24.84 ;
      RECT  46.93 28.62 47.38 29.07 ;
      RECT  48.77 24.37 48.91 26.68 ;
      RECT  47.89 25.71 48.03 29.29 ;
      RECT  48.68 26.68 49.03 27.03 ;
      RECT  47.89 33.55 48.03 32.56 ;
      RECT  48.77 30.89 48.91 28.63 ;
      RECT  47.89 32.56 48.24 32.21 ;
      RECT  46.93 33.53 47.38 33.08 ;
      RECT  46.93 29.3 47.38 28.85 ;
      RECT  48.77 33.55 48.91 31.24 ;
      RECT  47.89 32.21 48.03 28.63 ;
      RECT  48.68 31.24 49.03 30.89 ;
      RECT  47.89 33.07 48.03 34.06 ;
      RECT  48.77 35.73 48.91 37.99 ;
      RECT  47.89 34.06 48.24 34.41 ;
      RECT  46.93 33.09 47.38 33.54 ;
      RECT  46.93 37.32 47.38 37.77 ;
      RECT  48.77 33.07 48.91 35.38 ;
      RECT  47.89 34.41 48.03 37.99 ;
      RECT  48.68 35.38 49.03 35.73 ;
      RECT  47.89 42.25 48.03 41.26 ;
      RECT  48.77 39.59 48.91 37.33 ;
      RECT  47.89 41.26 48.24 40.91 ;
      RECT  46.93 42.23 47.38 41.78 ;
      RECT  46.93 38.0 47.38 37.55 ;
      RECT  48.77 42.25 48.91 39.94 ;
      RECT  47.89 40.91 48.03 37.33 ;
      RECT  48.68 39.94 49.03 39.59 ;
      RECT  47.89 41.77 48.03 42.76 ;
      RECT  48.77 44.43 48.91 46.69 ;
      RECT  47.89 42.76 48.24 43.11 ;
      RECT  46.93 41.79 47.38 42.24 ;
      RECT  46.93 46.02 47.38 46.47 ;
      RECT  48.77 41.77 48.91 44.08 ;
      RECT  47.89 43.11 48.03 46.69 ;
      RECT  48.68 44.08 49.03 44.43 ;
      RECT  47.89 50.95 48.03 49.96 ;
      RECT  48.77 48.29 48.91 46.03 ;
      RECT  47.89 49.96 48.24 49.61 ;
      RECT  46.93 50.93 47.38 50.48 ;
      RECT  46.93 46.7 47.38 46.25 ;
      RECT  48.77 50.95 48.91 48.64 ;
      RECT  47.89 49.61 48.03 46.03 ;
      RECT  48.68 48.64 49.03 48.29 ;
      RECT  47.89 50.47 48.03 51.46 ;
      RECT  48.77 53.13 48.91 55.39 ;
      RECT  47.89 51.46 48.24 51.81 ;
      RECT  46.93 50.49 47.38 50.94 ;
      RECT  46.93 54.72 47.38 55.17 ;
      RECT  48.77 50.47 48.91 52.78 ;
      RECT  47.89 51.81 48.03 55.39 ;
      RECT  48.68 52.78 49.03 53.13 ;
      RECT  47.89 59.65 48.03 58.66 ;
      RECT  48.77 56.99 48.91 54.73 ;
      RECT  47.89 58.66 48.24 58.31 ;
      RECT  46.93 59.63 47.38 59.18 ;
      RECT  46.93 55.4 47.38 54.95 ;
      RECT  48.77 59.65 48.91 57.34 ;
      RECT  47.89 58.31 48.03 54.73 ;
      RECT  48.68 57.34 49.03 56.99 ;
      RECT  47.89 59.17 48.03 60.16 ;
      RECT  48.77 61.83 48.91 64.09 ;
      RECT  47.89 60.16 48.24 60.51 ;
      RECT  46.93 59.19 47.38 59.64 ;
      RECT  46.93 63.42 47.38 63.87 ;
      RECT  48.77 59.17 48.91 61.48 ;
      RECT  47.89 60.51 48.03 64.09 ;
      RECT  48.68 61.48 49.03 61.83 ;
      RECT  47.89 68.35 48.03 67.36 ;
      RECT  48.77 65.69 48.91 63.43 ;
      RECT  47.89 67.36 48.24 67.01 ;
      RECT  46.93 68.33 47.38 67.88 ;
      RECT  46.93 64.1 47.38 63.65 ;
      RECT  48.77 68.35 48.91 66.04 ;
      RECT  47.89 67.01 48.03 63.43 ;
      RECT  48.68 66.04 49.03 65.69 ;
      RECT  47.89 67.87 48.03 68.86 ;
      RECT  48.77 70.53 48.91 72.79 ;
      RECT  47.89 68.86 48.24 69.21 ;
      RECT  46.93 67.89 47.38 68.34 ;
      RECT  46.93 72.12 47.38 72.57 ;
      RECT  48.77 67.87 48.91 70.18 ;
      RECT  47.89 69.21 48.03 72.79 ;
      RECT  48.68 70.18 49.03 70.53 ;
      RECT  47.89 77.05 48.03 76.06 ;
      RECT  48.77 74.39 48.91 72.13 ;
      RECT  47.89 76.06 48.24 75.71 ;
      RECT  46.93 77.03 47.38 76.58 ;
      RECT  46.93 72.8 47.38 72.35 ;
      RECT  48.77 77.05 48.91 74.74 ;
      RECT  47.89 75.71 48.03 72.13 ;
      RECT  48.68 74.74 49.03 74.39 ;
      RECT  47.89 76.57 48.03 77.56 ;
      RECT  48.77 79.23 48.91 81.49 ;
      RECT  47.89 77.56 48.24 77.91 ;
      RECT  46.93 76.59 47.38 77.04 ;
      RECT  46.93 80.82 47.38 81.27 ;
      RECT  48.77 76.57 48.91 78.88 ;
      RECT  47.89 77.91 48.03 81.49 ;
      RECT  48.68 78.88 49.03 79.23 ;
      RECT  47.89 85.75 48.03 84.76 ;
      RECT  48.77 83.09 48.91 80.83 ;
      RECT  47.89 84.76 48.24 84.41 ;
      RECT  46.93 85.73 47.38 85.28 ;
      RECT  46.93 81.5 47.38 81.05 ;
      RECT  48.77 85.75 48.91 83.44 ;
      RECT  47.89 84.41 48.03 80.83 ;
      RECT  48.68 83.44 49.03 83.09 ;
      RECT  47.89 85.27 48.03 86.26 ;
      RECT  48.77 87.93 48.91 90.19 ;
      RECT  47.89 86.26 48.24 86.61 ;
      RECT  46.93 85.29 47.38 85.74 ;
      RECT  46.93 89.52 47.38 89.97 ;
      RECT  48.77 85.27 48.91 87.58 ;
      RECT  47.89 86.61 48.03 90.19 ;
      RECT  48.68 87.58 49.03 87.93 ;
      RECT  47.89 94.45 48.03 93.46 ;
      RECT  48.77 91.79 48.91 89.53 ;
      RECT  47.89 93.46 48.24 93.11 ;
      RECT  46.93 94.43 47.38 93.98 ;
      RECT  46.93 90.2 47.38 89.75 ;
      RECT  48.77 94.45 48.91 92.14 ;
      RECT  47.89 93.11 48.03 89.53 ;
      RECT  48.68 92.14 49.03 91.79 ;
      RECT  47.89 93.97 48.03 94.96 ;
      RECT  48.77 96.63 48.91 98.89 ;
      RECT  47.89 94.96 48.24 95.31 ;
      RECT  46.93 93.99 47.38 94.44 ;
      RECT  46.93 98.22 47.38 98.67 ;
      RECT  48.77 93.97 48.91 96.28 ;
      RECT  47.89 95.31 48.03 98.89 ;
      RECT  48.68 96.28 49.03 96.63 ;
      RECT  47.89 103.15 48.03 102.16 ;
      RECT  48.77 100.49 48.91 98.23 ;
      RECT  47.89 102.16 48.24 101.81 ;
      RECT  46.93 103.13 47.38 102.68 ;
      RECT  46.93 98.9 47.38 98.45 ;
      RECT  48.77 103.15 48.91 100.84 ;
      RECT  47.89 101.81 48.03 98.23 ;
      RECT  48.68 100.84 49.03 100.49 ;
      RECT  47.89 102.67 48.03 103.66 ;
      RECT  48.77 105.33 48.91 107.59 ;
      RECT  47.89 103.66 48.24 104.01 ;
      RECT  46.93 102.69 47.38 103.14 ;
      RECT  46.93 106.92 47.38 107.37 ;
      RECT  48.77 102.67 48.91 104.98 ;
      RECT  47.89 104.01 48.03 107.59 ;
      RECT  48.68 104.98 49.03 105.33 ;
      RECT  47.89 24.61 48.24 107.26 ;
      RECT  48.68 24.61 49.03 107.26 ;
      RECT  50.97 33.55 51.11 32.56 ;
      RECT  51.85 30.89 51.99 28.63 ;
      RECT  50.97 32.56 51.32 32.21 ;
      RECT  50.01 33.53 50.46 33.08 ;
      RECT  50.01 29.3 50.46 28.85 ;
      RECT  51.85 33.55 51.99 31.24 ;
      RECT  50.97 32.21 51.11 28.63 ;
      RECT  51.76 31.24 52.11 30.89 ;
      RECT  54.05 33.55 54.19 32.56 ;
      RECT  54.93 30.89 55.07 28.63 ;
      RECT  54.05 32.56 54.4 32.21 ;
      RECT  53.09 33.53 53.54 33.08 ;
      RECT  53.09 29.3 53.54 28.85 ;
      RECT  54.93 33.55 55.07 31.24 ;
      RECT  54.05 32.21 54.19 28.63 ;
      RECT  54.84 31.24 55.19 30.89 ;
      RECT  50.97 33.31 51.32 28.96 ;
      RECT  51.76 33.31 52.11 28.96 ;
      RECT  54.05 33.31 54.4 28.96 ;
      RECT  54.84 33.31 55.19 28.96 ;
      RECT  50.97 24.37 51.11 25.36 ;
      RECT  51.85 27.03 51.99 29.29 ;
      RECT  50.97 25.36 51.32 25.71 ;
      RECT  50.01 24.39 50.46 24.84 ;
      RECT  50.01 28.62 50.46 29.07 ;
      RECT  51.85 24.37 51.99 26.68 ;
      RECT  50.97 25.71 51.11 29.29 ;
      RECT  51.76 26.68 52.11 27.03 ;
      RECT  54.05 24.37 54.19 25.36 ;
      RECT  54.93 27.03 55.07 29.29 ;
      RECT  54.05 25.36 54.4 25.71 ;
      RECT  53.09 24.39 53.54 24.84 ;
      RECT  53.09 28.62 53.54 29.07 ;
      RECT  54.93 24.37 55.07 26.68 ;
      RECT  54.05 25.71 54.19 29.29 ;
      RECT  54.84 26.68 55.19 27.03 ;
      RECT  50.97 24.61 51.32 28.96 ;
      RECT  51.76 24.61 52.11 28.96 ;
      RECT  54.05 24.61 54.4 28.96 ;
      RECT  54.84 24.61 55.19 28.96 ;
      RECT  50.97 102.67 51.11 103.66 ;
      RECT  51.85 105.33 51.99 107.59 ;
      RECT  50.97 103.66 51.32 104.01 ;
      RECT  50.01 102.69 50.46 103.14 ;
      RECT  50.01 106.92 50.46 107.37 ;
      RECT  51.85 102.67 51.99 104.98 ;
      RECT  50.97 104.01 51.11 107.59 ;
      RECT  51.76 104.98 52.11 105.33 ;
      RECT  54.05 102.67 54.19 103.66 ;
      RECT  54.93 105.33 55.07 107.59 ;
      RECT  54.05 103.66 54.4 104.01 ;
      RECT  53.09 102.69 53.54 103.14 ;
      RECT  53.09 106.92 53.54 107.37 ;
      RECT  54.93 102.67 55.07 104.98 ;
      RECT  54.05 104.01 54.19 107.59 ;
      RECT  54.84 104.98 55.19 105.33 ;
      RECT  50.97 102.91 51.32 107.26 ;
      RECT  51.76 102.91 52.11 107.26 ;
      RECT  54.05 102.91 54.4 107.26 ;
      RECT  54.84 102.91 55.19 107.26 ;
      RECT  44.81 24.37 44.95 25.36 ;
      RECT  45.69 27.03 45.83 29.29 ;
      RECT  44.81 25.36 45.16 25.71 ;
      RECT  43.85 24.39 44.3 24.84 ;
      RECT  43.85 28.62 44.3 29.07 ;
      RECT  45.69 24.37 45.83 26.68 ;
      RECT  44.81 25.71 44.95 29.29 ;
      RECT  45.6 26.68 45.95 27.03 ;
      RECT  44.81 33.55 44.95 32.56 ;
      RECT  45.69 30.89 45.83 28.63 ;
      RECT  44.81 32.56 45.16 32.21 ;
      RECT  43.85 33.53 44.3 33.08 ;
      RECT  43.85 29.3 44.3 28.85 ;
      RECT  45.69 33.55 45.83 31.24 ;
      RECT  44.81 32.21 44.95 28.63 ;
      RECT  45.6 31.24 45.95 30.89 ;
      RECT  44.81 33.07 44.95 34.06 ;
      RECT  45.69 35.73 45.83 37.99 ;
      RECT  44.81 34.06 45.16 34.41 ;
      RECT  43.85 33.09 44.3 33.54 ;
      RECT  43.85 37.32 44.3 37.77 ;
      RECT  45.69 33.07 45.83 35.38 ;
      RECT  44.81 34.41 44.95 37.99 ;
      RECT  45.6 35.38 45.95 35.73 ;
      RECT  44.81 42.25 44.95 41.26 ;
      RECT  45.69 39.59 45.83 37.33 ;
      RECT  44.81 41.26 45.16 40.91 ;
      RECT  43.85 42.23 44.3 41.78 ;
      RECT  43.85 38.0 44.3 37.55 ;
      RECT  45.69 42.25 45.83 39.94 ;
      RECT  44.81 40.91 44.95 37.33 ;
      RECT  45.6 39.94 45.95 39.59 ;
      RECT  44.81 41.77 44.95 42.76 ;
      RECT  45.69 44.43 45.83 46.69 ;
      RECT  44.81 42.76 45.16 43.11 ;
      RECT  43.85 41.79 44.3 42.24 ;
      RECT  43.85 46.02 44.3 46.47 ;
      RECT  45.69 41.77 45.83 44.08 ;
      RECT  44.81 43.11 44.95 46.69 ;
      RECT  45.6 44.08 45.95 44.43 ;
      RECT  44.81 50.95 44.95 49.96 ;
      RECT  45.69 48.29 45.83 46.03 ;
      RECT  44.81 49.96 45.16 49.61 ;
      RECT  43.85 50.93 44.3 50.48 ;
      RECT  43.85 46.7 44.3 46.25 ;
      RECT  45.69 50.95 45.83 48.64 ;
      RECT  44.81 49.61 44.95 46.03 ;
      RECT  45.6 48.64 45.95 48.29 ;
      RECT  44.81 50.47 44.95 51.46 ;
      RECT  45.69 53.13 45.83 55.39 ;
      RECT  44.81 51.46 45.16 51.81 ;
      RECT  43.85 50.49 44.3 50.94 ;
      RECT  43.85 54.72 44.3 55.17 ;
      RECT  45.69 50.47 45.83 52.78 ;
      RECT  44.81 51.81 44.95 55.39 ;
      RECT  45.6 52.78 45.95 53.13 ;
      RECT  44.81 59.65 44.95 58.66 ;
      RECT  45.69 56.99 45.83 54.73 ;
      RECT  44.81 58.66 45.16 58.31 ;
      RECT  43.85 59.63 44.3 59.18 ;
      RECT  43.85 55.4 44.3 54.95 ;
      RECT  45.69 59.65 45.83 57.34 ;
      RECT  44.81 58.31 44.95 54.73 ;
      RECT  45.6 57.34 45.95 56.99 ;
      RECT  44.81 59.17 44.95 60.16 ;
      RECT  45.69 61.83 45.83 64.09 ;
      RECT  44.81 60.16 45.16 60.51 ;
      RECT  43.85 59.19 44.3 59.64 ;
      RECT  43.85 63.42 44.3 63.87 ;
      RECT  45.69 59.17 45.83 61.48 ;
      RECT  44.81 60.51 44.95 64.09 ;
      RECT  45.6 61.48 45.95 61.83 ;
      RECT  44.81 68.35 44.95 67.36 ;
      RECT  45.69 65.69 45.83 63.43 ;
      RECT  44.81 67.36 45.16 67.01 ;
      RECT  43.85 68.33 44.3 67.88 ;
      RECT  43.85 64.1 44.3 63.65 ;
      RECT  45.69 68.35 45.83 66.04 ;
      RECT  44.81 67.01 44.95 63.43 ;
      RECT  45.6 66.04 45.95 65.69 ;
      RECT  44.81 67.87 44.95 68.86 ;
      RECT  45.69 70.53 45.83 72.79 ;
      RECT  44.81 68.86 45.16 69.21 ;
      RECT  43.85 67.89 44.3 68.34 ;
      RECT  43.85 72.12 44.3 72.57 ;
      RECT  45.69 67.87 45.83 70.18 ;
      RECT  44.81 69.21 44.95 72.79 ;
      RECT  45.6 70.18 45.95 70.53 ;
      RECT  44.81 77.05 44.95 76.06 ;
      RECT  45.69 74.39 45.83 72.13 ;
      RECT  44.81 76.06 45.16 75.71 ;
      RECT  43.85 77.03 44.3 76.58 ;
      RECT  43.85 72.8 44.3 72.35 ;
      RECT  45.69 77.05 45.83 74.74 ;
      RECT  44.81 75.71 44.95 72.13 ;
      RECT  45.6 74.74 45.95 74.39 ;
      RECT  44.81 76.57 44.95 77.56 ;
      RECT  45.69 79.23 45.83 81.49 ;
      RECT  44.81 77.56 45.16 77.91 ;
      RECT  43.85 76.59 44.3 77.04 ;
      RECT  43.85 80.82 44.3 81.27 ;
      RECT  45.69 76.57 45.83 78.88 ;
      RECT  44.81 77.91 44.95 81.49 ;
      RECT  45.6 78.88 45.95 79.23 ;
      RECT  44.81 85.75 44.95 84.76 ;
      RECT  45.69 83.09 45.83 80.83 ;
      RECT  44.81 84.76 45.16 84.41 ;
      RECT  43.85 85.73 44.3 85.28 ;
      RECT  43.85 81.5 44.3 81.05 ;
      RECT  45.69 85.75 45.83 83.44 ;
      RECT  44.81 84.41 44.95 80.83 ;
      RECT  45.6 83.44 45.95 83.09 ;
      RECT  44.81 85.27 44.95 86.26 ;
      RECT  45.69 87.93 45.83 90.19 ;
      RECT  44.81 86.26 45.16 86.61 ;
      RECT  43.85 85.29 44.3 85.74 ;
      RECT  43.85 89.52 44.3 89.97 ;
      RECT  45.69 85.27 45.83 87.58 ;
      RECT  44.81 86.61 44.95 90.19 ;
      RECT  45.6 87.58 45.95 87.93 ;
      RECT  44.81 94.45 44.95 93.46 ;
      RECT  45.69 91.79 45.83 89.53 ;
      RECT  44.81 93.46 45.16 93.11 ;
      RECT  43.85 94.43 44.3 93.98 ;
      RECT  43.85 90.2 44.3 89.75 ;
      RECT  45.69 94.45 45.83 92.14 ;
      RECT  44.81 93.11 44.95 89.53 ;
      RECT  45.6 92.14 45.95 91.79 ;
      RECT  44.81 93.97 44.95 94.96 ;
      RECT  45.69 96.63 45.83 98.89 ;
      RECT  44.81 94.96 45.16 95.31 ;
      RECT  43.85 93.99 44.3 94.44 ;
      RECT  43.85 98.22 44.3 98.67 ;
      RECT  45.69 93.97 45.83 96.28 ;
      RECT  44.81 95.31 44.95 98.89 ;
      RECT  45.6 96.28 45.95 96.63 ;
      RECT  44.81 103.15 44.95 102.16 ;
      RECT  45.69 100.49 45.83 98.23 ;
      RECT  44.81 102.16 45.16 101.81 ;
      RECT  43.85 103.13 44.3 102.68 ;
      RECT  43.85 98.9 44.3 98.45 ;
      RECT  45.69 103.15 45.83 100.84 ;
      RECT  44.81 101.81 44.95 98.23 ;
      RECT  45.6 100.84 45.95 100.49 ;
      RECT  44.81 102.67 44.95 103.66 ;
      RECT  45.69 105.33 45.83 107.59 ;
      RECT  44.81 103.66 45.16 104.01 ;
      RECT  43.85 102.69 44.3 103.14 ;
      RECT  43.85 106.92 44.3 107.37 ;
      RECT  45.69 102.67 45.83 104.98 ;
      RECT  44.81 104.01 44.95 107.59 ;
      RECT  45.6 104.98 45.95 105.33 ;
      RECT  44.81 24.61 45.16 107.26 ;
      RECT  45.6 24.61 45.95 107.26 ;
      RECT  57.13 24.37 57.27 25.36 ;
      RECT  58.01 27.03 58.15 29.29 ;
      RECT  57.13 25.36 57.48 25.71 ;
      RECT  56.17 24.39 56.62 24.84 ;
      RECT  56.17 28.62 56.62 29.07 ;
      RECT  58.01 24.37 58.15 26.68 ;
      RECT  57.13 25.71 57.27 29.29 ;
      RECT  57.92 26.68 58.27 27.03 ;
      RECT  57.13 33.55 57.27 32.56 ;
      RECT  58.01 30.89 58.15 28.63 ;
      RECT  57.13 32.56 57.48 32.21 ;
      RECT  56.17 33.53 56.62 33.08 ;
      RECT  56.17 29.3 56.62 28.85 ;
      RECT  58.01 33.55 58.15 31.24 ;
      RECT  57.13 32.21 57.27 28.63 ;
      RECT  57.92 31.24 58.27 30.89 ;
      RECT  57.13 33.07 57.27 34.06 ;
      RECT  58.01 35.73 58.15 37.99 ;
      RECT  57.13 34.06 57.48 34.41 ;
      RECT  56.17 33.09 56.62 33.54 ;
      RECT  56.17 37.32 56.62 37.77 ;
      RECT  58.01 33.07 58.15 35.38 ;
      RECT  57.13 34.41 57.27 37.99 ;
      RECT  57.92 35.38 58.27 35.73 ;
      RECT  57.13 42.25 57.27 41.26 ;
      RECT  58.01 39.59 58.15 37.33 ;
      RECT  57.13 41.26 57.48 40.91 ;
      RECT  56.17 42.23 56.62 41.78 ;
      RECT  56.17 38.0 56.62 37.55 ;
      RECT  58.01 42.25 58.15 39.94 ;
      RECT  57.13 40.91 57.27 37.33 ;
      RECT  57.92 39.94 58.27 39.59 ;
      RECT  57.13 41.77 57.27 42.76 ;
      RECT  58.01 44.43 58.15 46.69 ;
      RECT  57.13 42.76 57.48 43.11 ;
      RECT  56.17 41.79 56.62 42.24 ;
      RECT  56.17 46.02 56.62 46.47 ;
      RECT  58.01 41.77 58.15 44.08 ;
      RECT  57.13 43.11 57.27 46.69 ;
      RECT  57.92 44.08 58.27 44.43 ;
      RECT  57.13 50.95 57.27 49.96 ;
      RECT  58.01 48.29 58.15 46.03 ;
      RECT  57.13 49.96 57.48 49.61 ;
      RECT  56.17 50.93 56.62 50.48 ;
      RECT  56.17 46.7 56.62 46.25 ;
      RECT  58.01 50.95 58.15 48.64 ;
      RECT  57.13 49.61 57.27 46.03 ;
      RECT  57.92 48.64 58.27 48.29 ;
      RECT  57.13 50.47 57.27 51.46 ;
      RECT  58.01 53.13 58.15 55.39 ;
      RECT  57.13 51.46 57.48 51.81 ;
      RECT  56.17 50.49 56.62 50.94 ;
      RECT  56.17 54.72 56.62 55.17 ;
      RECT  58.01 50.47 58.15 52.78 ;
      RECT  57.13 51.81 57.27 55.39 ;
      RECT  57.92 52.78 58.27 53.13 ;
      RECT  57.13 59.65 57.27 58.66 ;
      RECT  58.01 56.99 58.15 54.73 ;
      RECT  57.13 58.66 57.48 58.31 ;
      RECT  56.17 59.63 56.62 59.18 ;
      RECT  56.17 55.4 56.62 54.95 ;
      RECT  58.01 59.65 58.15 57.34 ;
      RECT  57.13 58.31 57.27 54.73 ;
      RECT  57.92 57.34 58.27 56.99 ;
      RECT  57.13 59.17 57.27 60.16 ;
      RECT  58.01 61.83 58.15 64.09 ;
      RECT  57.13 60.16 57.48 60.51 ;
      RECT  56.17 59.19 56.62 59.64 ;
      RECT  56.17 63.42 56.62 63.87 ;
      RECT  58.01 59.17 58.15 61.48 ;
      RECT  57.13 60.51 57.27 64.09 ;
      RECT  57.92 61.48 58.27 61.83 ;
      RECT  57.13 68.35 57.27 67.36 ;
      RECT  58.01 65.69 58.15 63.43 ;
      RECT  57.13 67.36 57.48 67.01 ;
      RECT  56.17 68.33 56.62 67.88 ;
      RECT  56.17 64.1 56.62 63.65 ;
      RECT  58.01 68.35 58.15 66.04 ;
      RECT  57.13 67.01 57.27 63.43 ;
      RECT  57.92 66.04 58.27 65.69 ;
      RECT  57.13 67.87 57.27 68.86 ;
      RECT  58.01 70.53 58.15 72.79 ;
      RECT  57.13 68.86 57.48 69.21 ;
      RECT  56.17 67.89 56.62 68.34 ;
      RECT  56.17 72.12 56.62 72.57 ;
      RECT  58.01 67.87 58.15 70.18 ;
      RECT  57.13 69.21 57.27 72.79 ;
      RECT  57.92 70.18 58.27 70.53 ;
      RECT  57.13 77.05 57.27 76.06 ;
      RECT  58.01 74.39 58.15 72.13 ;
      RECT  57.13 76.06 57.48 75.71 ;
      RECT  56.17 77.03 56.62 76.58 ;
      RECT  56.17 72.8 56.62 72.35 ;
      RECT  58.01 77.05 58.15 74.74 ;
      RECT  57.13 75.71 57.27 72.13 ;
      RECT  57.92 74.74 58.27 74.39 ;
      RECT  57.13 76.57 57.27 77.56 ;
      RECT  58.01 79.23 58.15 81.49 ;
      RECT  57.13 77.56 57.48 77.91 ;
      RECT  56.17 76.59 56.62 77.04 ;
      RECT  56.17 80.82 56.62 81.27 ;
      RECT  58.01 76.57 58.15 78.88 ;
      RECT  57.13 77.91 57.27 81.49 ;
      RECT  57.92 78.88 58.27 79.23 ;
      RECT  57.13 85.75 57.27 84.76 ;
      RECT  58.01 83.09 58.15 80.83 ;
      RECT  57.13 84.76 57.48 84.41 ;
      RECT  56.17 85.73 56.62 85.28 ;
      RECT  56.17 81.5 56.62 81.05 ;
      RECT  58.01 85.75 58.15 83.44 ;
      RECT  57.13 84.41 57.27 80.83 ;
      RECT  57.92 83.44 58.27 83.09 ;
      RECT  57.13 85.27 57.27 86.26 ;
      RECT  58.01 87.93 58.15 90.19 ;
      RECT  57.13 86.26 57.48 86.61 ;
      RECT  56.17 85.29 56.62 85.74 ;
      RECT  56.17 89.52 56.62 89.97 ;
      RECT  58.01 85.27 58.15 87.58 ;
      RECT  57.13 86.61 57.27 90.19 ;
      RECT  57.92 87.58 58.27 87.93 ;
      RECT  57.13 94.45 57.27 93.46 ;
      RECT  58.01 91.79 58.15 89.53 ;
      RECT  57.13 93.46 57.48 93.11 ;
      RECT  56.17 94.43 56.62 93.98 ;
      RECT  56.17 90.2 56.62 89.75 ;
      RECT  58.01 94.45 58.15 92.14 ;
      RECT  57.13 93.11 57.27 89.53 ;
      RECT  57.92 92.14 58.27 91.79 ;
      RECT  57.13 93.97 57.27 94.96 ;
      RECT  58.01 96.63 58.15 98.89 ;
      RECT  57.13 94.96 57.48 95.31 ;
      RECT  56.17 93.99 56.62 94.44 ;
      RECT  56.17 98.22 56.62 98.67 ;
      RECT  58.01 93.97 58.15 96.28 ;
      RECT  57.13 95.31 57.27 98.89 ;
      RECT  57.92 96.28 58.27 96.63 ;
      RECT  57.13 103.15 57.27 102.16 ;
      RECT  58.01 100.49 58.15 98.23 ;
      RECT  57.13 102.16 57.48 101.81 ;
      RECT  56.17 103.13 56.62 102.68 ;
      RECT  56.17 98.9 56.62 98.45 ;
      RECT  58.01 103.15 58.15 100.84 ;
      RECT  57.13 101.81 57.27 98.23 ;
      RECT  57.92 100.84 58.27 100.49 ;
      RECT  57.13 102.67 57.27 103.66 ;
      RECT  58.01 105.33 58.15 107.59 ;
      RECT  57.13 103.66 57.48 104.01 ;
      RECT  56.17 102.69 56.62 103.14 ;
      RECT  56.17 106.92 56.62 107.37 ;
      RECT  58.01 102.67 58.15 104.98 ;
      RECT  57.13 104.01 57.27 107.59 ;
      RECT  57.92 104.98 58.27 105.33 ;
      RECT  57.13 24.61 57.48 107.26 ;
      RECT  57.92 24.61 58.27 107.26 ;
      RECT  47.89 24.61 48.24 107.26 ;
      RECT  48.68 24.61 49.03 107.26 ;
      RECT  50.97 24.61 51.32 107.26 ;
      RECT  51.76 24.61 52.11 107.26 ;
      RECT  54.05 24.61 54.4 107.26 ;
      RECT  54.84 24.61 55.19 107.26 ;
      RECT  47.12 15.63 47.26 22.63 ;
      RECT  48.88 15.63 49.02 22.63 ;
      RECT  50.2 15.63 50.34 22.63 ;
      RECT  51.96 15.63 52.1 22.63 ;
      RECT  53.28 15.63 53.42 22.63 ;
      RECT  55.04 15.63 55.18 22.63 ;
      RECT  47.12 15.63 47.26 22.63 ;
      RECT  48.88 15.63 49.02 22.63 ;
      RECT  50.2 15.63 50.34 22.63 ;
      RECT  51.96 15.63 52.1 22.63 ;
      RECT  53.28 15.63 53.42 22.63 ;
      RECT  55.04 15.63 55.18 22.63 ;
      RECT  49.84 13.42 50.29 13.87 ;
      RECT  49.96 8.83 50.41 9.28 ;
      RECT  50.86 10.61 51.21 10.96 ;
      RECT  50.95 10.96 51.12 14.09 ;
      RECT  52.2 11.02 52.55 11.37 ;
      RECT  52.29 11.37 52.46 14.09 ;
      RECT  50.95 8.81 51.12 10.61 ;
      RECT  52.29 8.81 52.46 11.02 ;
      RECT  52.92 13.42 53.37 13.87 ;
      RECT  53.04 8.83 53.49 9.28 ;
      RECT  53.94 10.61 54.29 10.96 ;
      RECT  54.03 10.96 54.2 14.09 ;
      RECT  55.28 11.02 55.63 11.37 ;
      RECT  55.37 11.37 55.54 14.09 ;
      RECT  54.03 8.81 54.2 10.61 ;
      RECT  55.37 8.81 55.54 11.02 ;
      RECT  50.86 10.61 51.21 10.96 ;
      RECT  52.2 11.02 52.55 11.37 ;
      RECT  53.94 10.61 54.29 10.96 ;
      RECT  55.28 11.02 55.63 11.37 ;
      RECT  51.39 -0.22 51.84 0.23 ;
      RECT  51.31 6.85 51.76 7.3 ;
      RECT  50.49 -0.25 50.77 1.45 ;
      RECT  52.13 1.31 52.41 7.33 ;
      RECT  49.89 1.8 50.04 6.48 ;
      RECT  52.13 -0.25 52.41 0.96 ;
      RECT  50.49 1.8 50.77 7.33 ;
      RECT  52.13 0.96 52.48 1.31 ;
      RECT  51.47 4.06 51.92 4.51 ;
      RECT  50.49 1.45 50.84 1.8 ;
      RECT  49.75 1.45 50.11 1.8 ;
      RECT  49.77 6.48 50.12 6.83 ;
      RECT  54.47 -0.22 54.92 0.23 ;
      RECT  54.39 6.85 54.84 7.3 ;
      RECT  53.57 -0.25 53.85 1.45 ;
      RECT  55.21 1.31 55.49 7.33 ;
      RECT  52.97 1.8 53.12 6.48 ;
      RECT  55.21 -0.25 55.49 0.96 ;
      RECT  53.57 1.8 53.85 7.33 ;
      RECT  55.21 0.96 55.56 1.31 ;
      RECT  54.55 4.06 55.0 4.51 ;
      RECT  53.57 1.45 53.92 1.8 ;
      RECT  52.83 1.45 53.19 1.8 ;
      RECT  52.85 6.48 53.2 6.83 ;
      RECT  50.49 1.45 50.84 1.8 ;
      RECT  52.13 0.96 52.48 1.31 ;
      RECT  53.57 1.45 53.92 1.8 ;
      RECT  55.21 0.96 55.56 1.31 ;
      RECT  47.12 22.63 47.26 15.63 ;
      RECT  48.88 22.63 49.02 15.63 ;
      RECT  50.2 22.63 50.34 15.63 ;
      RECT  51.96 22.63 52.1 15.63 ;
      RECT  53.28 22.63 53.42 15.63 ;
      RECT  55.04 22.63 55.18 15.63 ;
      RECT  3.44 35.15 3.9 35.61 ;
      RECT  4.1 39.71 4.56 40.17 ;
      RECT  3.44 61.25 3.9 61.71 ;
      RECT  4.1 65.81 4.56 66.27 ;
      RECT  0.16 33.31 0.3 76.81 ;
      RECT  0.82 33.31 0.96 76.81 ;
      RECT  1.48 33.31 1.62 76.81 ;
      RECT  2.14 33.31 2.28 76.81 ;
      RECT  34.585 33.31 34.725 102.91 ;
      RECT  0.16 33.31 0.3 76.81 ;
      RECT  0.82 33.31 0.96 76.81 ;
      RECT  1.48 33.31 1.62 76.81 ;
      RECT  2.14 33.31 2.28 76.81 ;
      RECT  34.09 31.725 34.23 31.865 ;
      RECT  0.16 33.31 0.3 76.81 ;
      RECT  0.82 33.31 0.96 76.81 ;
      RECT  1.48 33.31 1.62 76.81 ;
      RECT  2.14 33.31 2.28 76.81 ;
      RECT  37.63 0.0 37.77 24.61 ;
      RECT  39.27 0.0 39.41 24.61 ;
      RECT  38.45 0.0 38.59 24.61 ;
      RECT  40.09 0.0 40.23 24.61 ;
      RECT  -54.22 -6.98 -53.88 -6.66 ;
      RECT  -55.0 -7.8 -54.69 -7.48 ;
      RECT  -45.32 -7.29 -45.0 -6.97 ;
      RECT  -54.22 -6.98 -53.88 -6.66 ;
      RECT  -32.753 -8.795 -32.613 -8.655 ;
      RECT  -36.522 -6.12 -36.382 -5.98 ;
      RECT  -55.0 -7.8 -54.69 -7.48 ;
      RECT  -54.22 -3.46 -53.88 -3.78 ;
      RECT  -55.0 -2.64 -54.69 -2.96 ;
      RECT  -45.32 -3.15 -45.0 -3.47 ;
      RECT  -54.22 -3.46 -53.88 -3.78 ;
      RECT  -32.753 -1.645 -32.613 -1.785 ;
      RECT  -36.522 -4.32 -36.382 -4.46 ;
      RECT  -55.0 -2.64 -54.69 -2.96 ;
      RECT  -54.22 -6.98 -53.88 -6.66 ;
      RECT  -54.22 -3.78 -53.88 -3.46 ;
      RECT  -32.753 -8.795 -32.613 -8.655 ;
      RECT  -36.522 -6.12 -36.382 -5.98 ;
      RECT  -32.753 -1.785 -32.613 -1.645 ;
      RECT  -36.522 -4.46 -36.382 -4.32 ;
      RECT  -55.0 -9.31 -54.86 -1.13 ;
      RECT  -40.955 24.61 -41.095 28.705 ;
      RECT  -54.03 24.61 -54.17 95.905 ;
      RECT  -54.22 -6.98 -53.88 -6.66 ;
      RECT  -54.22 -3.78 -53.88 -3.46 ;
      RECT  -24.34 -7.44 -24.2 -7.3 ;
      RECT  -41.095 24.61 -40.955 28.705 ;
      RECT  -18.795 21.4 -1.32 21.54 ;
      RECT  -16.503 8.875 -1.32 9.015 ;
      RECT  -16.66 13.22 -1.32 13.36 ;
      RECT  -11.815 5.066 -1.32 5.206 ;
      RECT  -7.135 -7.493 -1.32 -7.353 ;
      RECT  -12.8 103.74 -12.46 104.06 ;
      RECT  -13.58 102.92 -13.27 103.24 ;
      RECT  -3.9 103.43 -3.58 103.75 ;
      RECT  -12.8 107.26 -12.46 106.94 ;
      RECT  -13.58 108.08 -13.27 107.76 ;
      RECT  -3.9 107.57 -3.58 107.25 ;
      RECT  -12.8 111.92 -12.46 112.24 ;
      RECT  -13.58 111.1 -13.27 111.42 ;
      RECT  -3.9 111.61 -3.58 111.93 ;
      RECT  -12.8 115.44 -12.46 115.12 ;
      RECT  -13.58 116.26 -13.27 115.94 ;
      RECT  -3.9 115.75 -3.58 115.43 ;
      RECT  -12.8 103.74 -12.46 104.06 ;
      RECT  -12.8 106.94 -12.46 107.26 ;
      RECT  -12.8 111.92 -12.46 112.24 ;
      RECT  -12.8 115.12 -12.46 115.44 ;
      RECT  -3.9 103.43 -3.58 103.75 ;
      RECT  -3.9 107.25 -3.58 107.57 ;
      RECT  -3.9 111.61 -3.58 111.93 ;
      RECT  -3.9 115.43 -3.58 115.75 ;
      RECT  12.62 -6.98 12.96 -6.66 ;
      RECT  11.84 -7.8 12.15 -7.48 ;
      RECT  21.52 -7.29 21.84 -6.97 ;
      RECT  25.33 -6.98 25.67 -6.66 ;
      RECT  24.55 -7.8 24.86 -7.48 ;
      RECT  34.23 -7.29 34.55 -6.97 ;
      RECT  12.62 -6.98 12.96 -6.66 ;
      RECT  25.33 -6.98 25.67 -6.66 ;
      RECT  21.52 -7.29 21.84 -6.97 ;
      RECT  34.23 -7.29 34.55 -6.97 ;
   LAYER  m3 ;
      RECT  49.99 33.07 50.47 33.16 ;
      RECT  49.61 33.16 52.69 33.46 ;
      RECT  49.99 33.46 50.48 33.56 ;
      RECT  49.97 37.28 50.5 37.51 ;
      RECT  49.61 37.51 52.69 37.81 ;
      RECT  49.99 42.25 50.47 42.16 ;
      RECT  49.61 42.16 52.69 41.86 ;
      RECT  49.99 41.86 50.48 41.76 ;
      RECT  49.97 38.04 50.5 37.81 ;
      RECT  49.61 37.81 52.69 37.51 ;
      RECT  49.99 41.77 50.47 41.86 ;
      RECT  49.61 41.86 52.69 42.16 ;
      RECT  49.99 42.16 50.48 42.26 ;
      RECT  49.97 45.98 50.5 46.21 ;
      RECT  49.61 46.21 52.69 46.51 ;
      RECT  49.99 50.95 50.47 50.86 ;
      RECT  49.61 50.86 52.69 50.56 ;
      RECT  49.99 50.56 50.48 50.46 ;
      RECT  49.97 46.74 50.5 46.51 ;
      RECT  49.61 46.51 52.69 46.21 ;
      RECT  49.99 50.47 50.47 50.56 ;
      RECT  49.61 50.56 52.69 50.86 ;
      RECT  49.99 50.86 50.48 50.96 ;
      RECT  49.97 54.68 50.5 54.91 ;
      RECT  49.61 54.91 52.69 55.21 ;
      RECT  49.99 59.65 50.47 59.56 ;
      RECT  49.61 59.56 52.69 59.26 ;
      RECT  49.99 59.26 50.48 59.16 ;
      RECT  49.97 55.44 50.5 55.21 ;
      RECT  49.61 55.21 52.69 54.91 ;
      RECT  49.99 59.17 50.47 59.26 ;
      RECT  49.61 59.26 52.69 59.56 ;
      RECT  49.99 59.56 50.48 59.66 ;
      RECT  49.97 63.38 50.5 63.61 ;
      RECT  49.61 63.61 52.69 63.91 ;
      RECT  49.99 68.35 50.47 68.26 ;
      RECT  49.61 68.26 52.69 67.96 ;
      RECT  49.99 67.96 50.48 67.86 ;
      RECT  49.97 64.14 50.5 63.91 ;
      RECT  49.61 63.91 52.69 63.61 ;
      RECT  49.99 67.87 50.47 67.96 ;
      RECT  49.61 67.96 52.69 68.26 ;
      RECT  49.99 68.26 50.48 68.36 ;
      RECT  49.97 72.08 50.5 72.31 ;
      RECT  49.61 72.31 52.69 72.61 ;
      RECT  49.99 77.05 50.47 76.96 ;
      RECT  49.61 76.96 52.69 76.66 ;
      RECT  49.99 76.66 50.48 76.56 ;
      RECT  49.97 72.84 50.5 72.61 ;
      RECT  49.61 72.61 52.69 72.31 ;
      RECT  49.99 76.57 50.47 76.66 ;
      RECT  49.61 76.66 52.69 76.96 ;
      RECT  49.99 76.96 50.48 77.06 ;
      RECT  49.97 80.78 50.5 81.01 ;
      RECT  49.61 81.01 52.69 81.31 ;
      RECT  49.99 85.75 50.47 85.66 ;
      RECT  49.61 85.66 52.69 85.36 ;
      RECT  49.99 85.36 50.48 85.26 ;
      RECT  49.97 81.54 50.5 81.31 ;
      RECT  49.61 81.31 52.69 81.01 ;
      RECT  49.99 85.27 50.47 85.36 ;
      RECT  49.61 85.36 52.69 85.66 ;
      RECT  49.99 85.66 50.48 85.76 ;
      RECT  49.97 89.48 50.5 89.71 ;
      RECT  49.61 89.71 52.69 90.01 ;
      RECT  49.99 94.45 50.47 94.36 ;
      RECT  49.61 94.36 52.69 94.06 ;
      RECT  49.99 94.06 50.48 93.96 ;
      RECT  49.97 90.24 50.5 90.01 ;
      RECT  49.61 90.01 52.69 89.71 ;
      RECT  49.99 93.97 50.47 94.06 ;
      RECT  49.61 94.06 52.69 94.36 ;
      RECT  49.99 94.36 50.48 94.46 ;
      RECT  49.97 98.18 50.5 98.41 ;
      RECT  49.61 98.41 52.69 98.71 ;
      RECT  49.99 103.15 50.47 103.06 ;
      RECT  49.61 103.06 52.69 102.76 ;
      RECT  49.99 102.76 50.48 102.66 ;
      RECT  49.97 98.94 50.5 98.71 ;
      RECT  49.61 98.71 52.69 98.41 ;
      RECT  53.07 33.07 53.55 33.16 ;
      RECT  52.69 33.16 55.77 33.46 ;
      RECT  53.07 33.46 53.56 33.56 ;
      RECT  53.05 37.28 53.58 37.51 ;
      RECT  52.69 37.51 55.77 37.81 ;
      RECT  53.07 42.25 53.55 42.16 ;
      RECT  52.69 42.16 55.77 41.86 ;
      RECT  53.07 41.86 53.56 41.76 ;
      RECT  53.05 38.04 53.58 37.81 ;
      RECT  52.69 37.81 55.77 37.51 ;
      RECT  53.07 41.77 53.55 41.86 ;
      RECT  52.69 41.86 55.77 42.16 ;
      RECT  53.07 42.16 53.56 42.26 ;
      RECT  53.05 45.98 53.58 46.21 ;
      RECT  52.69 46.21 55.77 46.51 ;
      RECT  53.07 50.95 53.55 50.86 ;
      RECT  52.69 50.86 55.77 50.56 ;
      RECT  53.07 50.56 53.56 50.46 ;
      RECT  53.05 46.74 53.58 46.51 ;
      RECT  52.69 46.51 55.77 46.21 ;
      RECT  53.07 50.47 53.55 50.56 ;
      RECT  52.69 50.56 55.77 50.86 ;
      RECT  53.07 50.86 53.56 50.96 ;
      RECT  53.05 54.68 53.58 54.91 ;
      RECT  52.69 54.91 55.77 55.21 ;
      RECT  53.07 59.65 53.55 59.56 ;
      RECT  52.69 59.56 55.77 59.26 ;
      RECT  53.07 59.26 53.56 59.16 ;
      RECT  53.05 55.44 53.58 55.21 ;
      RECT  52.69 55.21 55.77 54.91 ;
      RECT  53.07 59.17 53.55 59.26 ;
      RECT  52.69 59.26 55.77 59.56 ;
      RECT  53.07 59.56 53.56 59.66 ;
      RECT  53.05 63.38 53.58 63.61 ;
      RECT  52.69 63.61 55.77 63.91 ;
      RECT  53.07 68.35 53.55 68.26 ;
      RECT  52.69 68.26 55.77 67.96 ;
      RECT  53.07 67.96 53.56 67.86 ;
      RECT  53.05 64.14 53.58 63.91 ;
      RECT  52.69 63.91 55.77 63.61 ;
      RECT  53.07 67.87 53.55 67.96 ;
      RECT  52.69 67.96 55.77 68.26 ;
      RECT  53.07 68.26 53.56 68.36 ;
      RECT  53.05 72.08 53.58 72.31 ;
      RECT  52.69 72.31 55.77 72.61 ;
      RECT  53.07 77.05 53.55 76.96 ;
      RECT  52.69 76.96 55.77 76.66 ;
      RECT  53.07 76.66 53.56 76.56 ;
      RECT  53.05 72.84 53.58 72.61 ;
      RECT  52.69 72.61 55.77 72.31 ;
      RECT  53.07 76.57 53.55 76.66 ;
      RECT  52.69 76.66 55.77 76.96 ;
      RECT  53.07 76.96 53.56 77.06 ;
      RECT  53.05 80.78 53.58 81.01 ;
      RECT  52.69 81.01 55.77 81.31 ;
      RECT  53.07 85.75 53.55 85.66 ;
      RECT  52.69 85.66 55.77 85.36 ;
      RECT  53.07 85.36 53.56 85.26 ;
      RECT  53.05 81.54 53.58 81.31 ;
      RECT  52.69 81.31 55.77 81.01 ;
      RECT  53.07 85.27 53.55 85.36 ;
      RECT  52.69 85.36 55.77 85.66 ;
      RECT  53.07 85.66 53.56 85.76 ;
      RECT  53.05 89.48 53.58 89.71 ;
      RECT  52.69 89.71 55.77 90.01 ;
      RECT  53.07 94.45 53.55 94.36 ;
      RECT  52.69 94.36 55.77 94.06 ;
      RECT  53.07 94.06 53.56 93.96 ;
      RECT  53.05 90.24 53.58 90.01 ;
      RECT  52.69 90.01 55.77 89.71 ;
      RECT  53.07 93.97 53.55 94.06 ;
      RECT  52.69 94.06 55.77 94.36 ;
      RECT  53.07 94.36 53.56 94.46 ;
      RECT  53.05 98.18 53.58 98.41 ;
      RECT  52.69 98.41 55.77 98.71 ;
      RECT  53.07 103.15 53.55 103.06 ;
      RECT  52.69 103.06 55.77 102.76 ;
      RECT  53.07 102.76 53.56 102.66 ;
      RECT  53.05 98.94 53.58 98.71 ;
      RECT  52.69 98.71 55.77 98.41 ;
      RECT  49.61 72.31 52.69 72.61 ;
      RECT  49.61 46.21 52.69 46.51 ;
      RECT  49.61 46.21 52.69 46.51 ;
      RECT  49.61 81.01 52.69 81.31 ;
      RECT  49.61 89.71 52.69 90.01 ;
      RECT  52.69 46.21 55.77 46.51 ;
      RECT  52.69 46.21 55.77 46.51 ;
      RECT  49.61 89.71 52.69 90.01 ;
      RECT  52.69 98.41 55.77 98.71 ;
      RECT  52.69 72.31 55.77 72.61 ;
      RECT  52.69 72.31 55.77 72.61 ;
      RECT  49.61 54.91 52.69 55.21 ;
      RECT  49.61 37.51 52.69 37.81 ;
      RECT  49.61 37.51 52.69 37.81 ;
      RECT  52.69 89.71 55.77 90.01 ;
      RECT  52.69 89.71 55.77 90.01 ;
      RECT  52.69 54.91 55.77 55.21 ;
      RECT  49.61 63.61 52.69 63.91 ;
      RECT  49.61 98.41 52.69 98.71 ;
      RECT  52.69 37.51 55.77 37.81 ;
      RECT  52.69 37.51 55.77 37.81 ;
      RECT  49.61 98.41 52.69 98.71 ;
      RECT  52.69 63.61 55.77 63.91 ;
      RECT  52.69 63.61 55.77 63.91 ;
      RECT  52.69 81.01 55.77 81.31 ;
      RECT  49.61 72.31 52.69 72.61 ;
      RECT  49.61 63.61 52.69 63.91 ;
      RECT  52.69 98.41 55.77 98.71 ;
      RECT  49.61 94.06 52.69 94.36 ;
      RECT  49.61 50.56 52.69 50.86 ;
      RECT  49.61 41.86 52.69 42.16 ;
      RECT  52.69 94.06 55.77 94.36 ;
      RECT  52.69 102.76 55.77 103.06 ;
      RECT  52.69 33.16 55.77 33.46 ;
      RECT  52.69 50.56 55.77 50.86 ;
      RECT  49.61 59.26 52.69 59.56 ;
      RECT  52.69 67.96 55.77 68.26 ;
      RECT  49.61 85.36 52.69 85.66 ;
      RECT  52.69 76.66 55.77 76.96 ;
      RECT  49.61 33.16 52.69 33.46 ;
      RECT  49.61 102.76 52.69 103.06 ;
      RECT  52.69 41.86 55.77 42.16 ;
      RECT  49.61 67.96 52.69 68.26 ;
      RECT  52.69 59.26 55.77 59.56 ;
      RECT  52.69 85.36 55.77 85.66 ;
      RECT  49.61 76.66 52.69 76.96 ;
      RECT  46.91 24.37 47.39 24.46 ;
      RECT  46.53 24.46 49.61 24.76 ;
      RECT  46.91 24.76 47.4 24.86 ;
      RECT  46.89 28.58 47.42 28.81 ;
      RECT  46.53 28.81 49.61 29.11 ;
      RECT  46.91 33.55 47.39 33.46 ;
      RECT  46.53 33.46 49.61 33.16 ;
      RECT  46.91 33.16 47.4 33.06 ;
      RECT  46.89 29.34 47.42 29.11 ;
      RECT  46.53 29.11 49.61 28.81 ;
      RECT  46.91 33.07 47.39 33.16 ;
      RECT  46.53 33.16 49.61 33.46 ;
      RECT  46.91 33.46 47.4 33.56 ;
      RECT  46.89 37.28 47.42 37.51 ;
      RECT  46.53 37.51 49.61 37.81 ;
      RECT  46.91 42.25 47.39 42.16 ;
      RECT  46.53 42.16 49.61 41.86 ;
      RECT  46.91 41.86 47.4 41.76 ;
      RECT  46.89 38.04 47.42 37.81 ;
      RECT  46.53 37.81 49.61 37.51 ;
      RECT  46.91 41.77 47.39 41.86 ;
      RECT  46.53 41.86 49.61 42.16 ;
      RECT  46.91 42.16 47.4 42.26 ;
      RECT  46.89 45.98 47.42 46.21 ;
      RECT  46.53 46.21 49.61 46.51 ;
      RECT  46.91 50.95 47.39 50.86 ;
      RECT  46.53 50.86 49.61 50.56 ;
      RECT  46.91 50.56 47.4 50.46 ;
      RECT  46.89 46.74 47.42 46.51 ;
      RECT  46.53 46.51 49.61 46.21 ;
      RECT  46.91 50.47 47.39 50.56 ;
      RECT  46.53 50.56 49.61 50.86 ;
      RECT  46.91 50.86 47.4 50.96 ;
      RECT  46.89 54.68 47.42 54.91 ;
      RECT  46.53 54.91 49.61 55.21 ;
      RECT  46.91 59.65 47.39 59.56 ;
      RECT  46.53 59.56 49.61 59.26 ;
      RECT  46.91 59.26 47.4 59.16 ;
      RECT  46.89 55.44 47.42 55.21 ;
      RECT  46.53 55.21 49.61 54.91 ;
      RECT  46.91 59.17 47.39 59.26 ;
      RECT  46.53 59.26 49.61 59.56 ;
      RECT  46.91 59.56 47.4 59.66 ;
      RECT  46.89 63.38 47.42 63.61 ;
      RECT  46.53 63.61 49.61 63.91 ;
      RECT  46.91 68.35 47.39 68.26 ;
      RECT  46.53 68.26 49.61 67.96 ;
      RECT  46.91 67.96 47.4 67.86 ;
      RECT  46.89 64.14 47.42 63.91 ;
      RECT  46.53 63.91 49.61 63.61 ;
      RECT  46.91 67.87 47.39 67.96 ;
      RECT  46.53 67.96 49.61 68.26 ;
      RECT  46.91 68.26 47.4 68.36 ;
      RECT  46.89 72.08 47.42 72.31 ;
      RECT  46.53 72.31 49.61 72.61 ;
      RECT  46.91 77.05 47.39 76.96 ;
      RECT  46.53 76.96 49.61 76.66 ;
      RECT  46.91 76.66 47.4 76.56 ;
      RECT  46.89 72.84 47.42 72.61 ;
      RECT  46.53 72.61 49.61 72.31 ;
      RECT  46.91 76.57 47.39 76.66 ;
      RECT  46.53 76.66 49.61 76.96 ;
      RECT  46.91 76.96 47.4 77.06 ;
      RECT  46.89 80.78 47.42 81.01 ;
      RECT  46.53 81.01 49.61 81.31 ;
      RECT  46.91 85.75 47.39 85.66 ;
      RECT  46.53 85.66 49.61 85.36 ;
      RECT  46.91 85.36 47.4 85.26 ;
      RECT  46.89 81.54 47.42 81.31 ;
      RECT  46.53 81.31 49.61 81.01 ;
      RECT  46.91 85.27 47.39 85.36 ;
      RECT  46.53 85.36 49.61 85.66 ;
      RECT  46.91 85.66 47.4 85.76 ;
      RECT  46.89 89.48 47.42 89.71 ;
      RECT  46.53 89.71 49.61 90.01 ;
      RECT  46.91 94.45 47.39 94.36 ;
      RECT  46.53 94.36 49.61 94.06 ;
      RECT  46.91 94.06 47.4 93.96 ;
      RECT  46.89 90.24 47.42 90.01 ;
      RECT  46.53 90.01 49.61 89.71 ;
      RECT  46.91 93.97 47.39 94.06 ;
      RECT  46.53 94.06 49.61 94.36 ;
      RECT  46.91 94.36 47.4 94.46 ;
      RECT  46.89 98.18 47.42 98.41 ;
      RECT  46.53 98.41 49.61 98.71 ;
      RECT  46.91 103.15 47.39 103.06 ;
      RECT  46.53 103.06 49.61 102.76 ;
      RECT  46.91 102.76 47.4 102.66 ;
      RECT  46.89 98.94 47.42 98.71 ;
      RECT  46.53 98.71 49.61 98.41 ;
      RECT  46.91 102.67 47.39 102.76 ;
      RECT  46.53 102.76 49.61 103.06 ;
      RECT  46.91 103.06 47.4 103.16 ;
      RECT  46.89 106.88 47.42 107.11 ;
      RECT  46.53 107.11 49.61 107.41 ;
      RECT  46.53 98.41 49.61 98.71 ;
      RECT  46.53 98.41 49.61 98.71 ;
      RECT  46.53 54.91 49.61 55.21 ;
      RECT  46.53 46.21 49.61 46.51 ;
      RECT  47.92 107.11 48.22 107.41 ;
      RECT  47.92 28.81 48.22 29.11 ;
      RECT  46.53 63.61 49.61 63.91 ;
      RECT  46.53 37.51 49.61 37.81 ;
      RECT  46.53 37.51 49.61 37.81 ;
      RECT  46.53 28.81 49.61 29.11 ;
      RECT  46.53 72.31 49.61 72.61 ;
      RECT  46.53 81.01 49.61 81.31 ;
      RECT  46.53 81.01 49.61 81.31 ;
      RECT  46.53 89.71 49.61 90.01 ;
      RECT  46.53 63.61 49.61 63.91 ;
      RECT  46.53 89.71 49.61 90.01 ;
      RECT  46.53 54.91 49.61 55.21 ;
      RECT  46.53 85.36 49.61 85.66 ;
      RECT  46.53 41.86 49.61 42.16 ;
      RECT  46.53 33.16 49.61 33.46 ;
      RECT  47.92 102.76 48.22 103.06 ;
      RECT  46.53 50.56 49.61 50.86 ;
      RECT  46.53 76.66 49.61 76.96 ;
      RECT  46.53 94.06 49.61 94.36 ;
      RECT  46.53 59.26 49.61 59.56 ;
      RECT  47.92 24.46 48.22 24.76 ;
      RECT  46.53 102.76 49.61 103.06 ;
      RECT  46.53 67.96 49.61 68.26 ;
      RECT  49.99 33.55 50.47 33.46 ;
      RECT  49.61 33.46 52.69 33.16 ;
      RECT  49.99 33.16 50.48 33.06 ;
      RECT  49.97 29.34 50.5 29.11 ;
      RECT  49.61 29.11 52.69 28.81 ;
      RECT  53.07 33.55 53.55 33.46 ;
      RECT  52.69 33.46 55.77 33.16 ;
      RECT  53.07 33.16 53.56 33.06 ;
      RECT  53.05 29.34 53.58 29.11 ;
      RECT  52.69 29.11 55.77 28.81 ;
      RECT  52.69 29.11 55.77 28.81 ;
      RECT  49.61 29.11 52.69 28.81 ;
      RECT  49.61 33.46 52.69 33.16 ;
      RECT  52.69 33.46 55.77 33.16 ;
      RECT  49.99 24.37 50.47 24.46 ;
      RECT  49.61 24.46 52.69 24.76 ;
      RECT  49.99 24.76 50.48 24.86 ;
      RECT  49.97 28.58 50.5 28.81 ;
      RECT  49.61 28.81 52.69 29.11 ;
      RECT  53.07 24.37 53.55 24.46 ;
      RECT  52.69 24.46 55.77 24.76 ;
      RECT  53.07 24.76 53.56 24.86 ;
      RECT  53.05 28.58 53.58 28.81 ;
      RECT  52.69 28.81 55.77 29.11 ;
      RECT  52.69 28.81 55.77 29.11 ;
      RECT  49.61 28.81 52.69 29.11 ;
      RECT  49.61 24.46 52.69 24.76 ;
      RECT  52.69 24.46 55.77 24.76 ;
      RECT  49.99 102.67 50.47 102.76 ;
      RECT  49.61 102.76 52.69 103.06 ;
      RECT  49.99 103.06 50.48 103.16 ;
      RECT  49.97 106.88 50.5 107.11 ;
      RECT  49.61 107.11 52.69 107.41 ;
      RECT  53.07 102.67 53.55 102.76 ;
      RECT  52.69 102.76 55.77 103.06 ;
      RECT  53.07 103.06 53.56 103.16 ;
      RECT  53.05 106.88 53.58 107.11 ;
      RECT  52.69 107.11 55.77 107.41 ;
      RECT  52.69 107.11 55.77 107.41 ;
      RECT  49.61 107.11 52.69 107.41 ;
      RECT  49.61 102.76 52.69 103.06 ;
      RECT  52.69 102.76 55.77 103.06 ;
      RECT  43.83 24.37 44.31 24.46 ;
      RECT  43.45 24.46 46.53 24.76 ;
      RECT  43.83 24.76 44.32 24.86 ;
      RECT  43.81 28.58 44.34 28.81 ;
      RECT  43.45 28.81 46.53 29.11 ;
      RECT  43.83 33.55 44.31 33.46 ;
      RECT  43.45 33.46 46.53 33.16 ;
      RECT  43.83 33.16 44.32 33.06 ;
      RECT  43.81 29.34 44.34 29.11 ;
      RECT  43.45 29.11 46.53 28.81 ;
      RECT  43.83 33.07 44.31 33.16 ;
      RECT  43.45 33.16 46.53 33.46 ;
      RECT  43.83 33.46 44.32 33.56 ;
      RECT  43.81 37.28 44.34 37.51 ;
      RECT  43.45 37.51 46.53 37.81 ;
      RECT  43.83 42.25 44.31 42.16 ;
      RECT  43.45 42.16 46.53 41.86 ;
      RECT  43.83 41.86 44.32 41.76 ;
      RECT  43.81 38.04 44.34 37.81 ;
      RECT  43.45 37.81 46.53 37.51 ;
      RECT  43.83 41.77 44.31 41.86 ;
      RECT  43.45 41.86 46.53 42.16 ;
      RECT  43.83 42.16 44.32 42.26 ;
      RECT  43.81 45.98 44.34 46.21 ;
      RECT  43.45 46.21 46.53 46.51 ;
      RECT  43.83 50.95 44.31 50.86 ;
      RECT  43.45 50.86 46.53 50.56 ;
      RECT  43.83 50.56 44.32 50.46 ;
      RECT  43.81 46.74 44.34 46.51 ;
      RECT  43.45 46.51 46.53 46.21 ;
      RECT  43.83 50.47 44.31 50.56 ;
      RECT  43.45 50.56 46.53 50.86 ;
      RECT  43.83 50.86 44.32 50.96 ;
      RECT  43.81 54.68 44.34 54.91 ;
      RECT  43.45 54.91 46.53 55.21 ;
      RECT  43.83 59.65 44.31 59.56 ;
      RECT  43.45 59.56 46.53 59.26 ;
      RECT  43.83 59.26 44.32 59.16 ;
      RECT  43.81 55.44 44.34 55.21 ;
      RECT  43.45 55.21 46.53 54.91 ;
      RECT  43.83 59.17 44.31 59.26 ;
      RECT  43.45 59.26 46.53 59.56 ;
      RECT  43.83 59.56 44.32 59.66 ;
      RECT  43.81 63.38 44.34 63.61 ;
      RECT  43.45 63.61 46.53 63.91 ;
      RECT  43.83 68.35 44.31 68.26 ;
      RECT  43.45 68.26 46.53 67.96 ;
      RECT  43.83 67.96 44.32 67.86 ;
      RECT  43.81 64.14 44.34 63.91 ;
      RECT  43.45 63.91 46.53 63.61 ;
      RECT  43.83 67.87 44.31 67.96 ;
      RECT  43.45 67.96 46.53 68.26 ;
      RECT  43.83 68.26 44.32 68.36 ;
      RECT  43.81 72.08 44.34 72.31 ;
      RECT  43.45 72.31 46.53 72.61 ;
      RECT  43.83 77.05 44.31 76.96 ;
      RECT  43.45 76.96 46.53 76.66 ;
      RECT  43.83 76.66 44.32 76.56 ;
      RECT  43.81 72.84 44.34 72.61 ;
      RECT  43.45 72.61 46.53 72.31 ;
      RECT  43.83 76.57 44.31 76.66 ;
      RECT  43.45 76.66 46.53 76.96 ;
      RECT  43.83 76.96 44.32 77.06 ;
      RECT  43.81 80.78 44.34 81.01 ;
      RECT  43.45 81.01 46.53 81.31 ;
      RECT  43.83 85.75 44.31 85.66 ;
      RECT  43.45 85.66 46.53 85.36 ;
      RECT  43.83 85.36 44.32 85.26 ;
      RECT  43.81 81.54 44.34 81.31 ;
      RECT  43.45 81.31 46.53 81.01 ;
      RECT  43.83 85.27 44.31 85.36 ;
      RECT  43.45 85.36 46.53 85.66 ;
      RECT  43.83 85.66 44.32 85.76 ;
      RECT  43.81 89.48 44.34 89.71 ;
      RECT  43.45 89.71 46.53 90.01 ;
      RECT  43.83 94.45 44.31 94.36 ;
      RECT  43.45 94.36 46.53 94.06 ;
      RECT  43.83 94.06 44.32 93.96 ;
      RECT  43.81 90.24 44.34 90.01 ;
      RECT  43.45 90.01 46.53 89.71 ;
      RECT  43.83 93.97 44.31 94.06 ;
      RECT  43.45 94.06 46.53 94.36 ;
      RECT  43.83 94.36 44.32 94.46 ;
      RECT  43.81 98.18 44.34 98.41 ;
      RECT  43.45 98.41 46.53 98.71 ;
      RECT  43.83 103.15 44.31 103.06 ;
      RECT  43.45 103.06 46.53 102.76 ;
      RECT  43.83 102.76 44.32 102.66 ;
      RECT  43.81 98.94 44.34 98.71 ;
      RECT  43.45 98.71 46.53 98.41 ;
      RECT  43.83 102.67 44.31 102.76 ;
      RECT  43.45 102.76 46.53 103.06 ;
      RECT  43.83 103.06 44.32 103.16 ;
      RECT  43.81 106.88 44.34 107.11 ;
      RECT  43.45 107.11 46.53 107.41 ;
      RECT  43.45 98.41 46.53 98.71 ;
      RECT  43.45 98.41 46.53 98.71 ;
      RECT  43.45 54.91 46.53 55.21 ;
      RECT  43.45 46.21 46.53 46.51 ;
      RECT  43.45 63.61 46.53 63.91 ;
      RECT  43.45 37.51 46.53 37.81 ;
      RECT  43.45 37.51 46.53 37.81 ;
      RECT  43.45 28.81 46.53 29.11 ;
      RECT  43.45 28.81 46.53 29.11 ;
      RECT  43.45 72.31 46.53 72.61 ;
      RECT  43.45 81.01 46.53 81.31 ;
      RECT  43.45 81.01 46.53 81.31 ;
      RECT  43.45 107.11 46.53 107.41 ;
      RECT  43.45 89.71 46.53 90.01 ;
      RECT  43.45 63.61 46.53 63.91 ;
      RECT  43.45 89.71 46.53 90.01 ;
      RECT  43.45 54.91 46.53 55.21 ;
      RECT  43.45 85.36 46.53 85.66 ;
      RECT  43.45 41.86 46.53 42.16 ;
      RECT  43.45 33.16 46.53 33.46 ;
      RECT  43.45 50.56 46.53 50.86 ;
      RECT  43.45 76.66 46.53 76.96 ;
      RECT  43.45 24.46 46.53 24.76 ;
      RECT  43.45 94.06 46.53 94.36 ;
      RECT  43.45 59.26 46.53 59.56 ;
      RECT  43.45 102.76 46.53 103.06 ;
      RECT  43.45 67.96 46.53 68.26 ;
      RECT  56.15 24.37 56.63 24.46 ;
      RECT  55.77 24.46 58.85 24.76 ;
      RECT  56.15 24.76 56.64 24.86 ;
      RECT  56.13 28.58 56.66 28.81 ;
      RECT  55.77 28.81 58.85 29.11 ;
      RECT  56.15 33.55 56.63 33.46 ;
      RECT  55.77 33.46 58.85 33.16 ;
      RECT  56.15 33.16 56.64 33.06 ;
      RECT  56.13 29.34 56.66 29.11 ;
      RECT  55.77 29.11 58.85 28.81 ;
      RECT  56.15 33.07 56.63 33.16 ;
      RECT  55.77 33.16 58.85 33.46 ;
      RECT  56.15 33.46 56.64 33.56 ;
      RECT  56.13 37.28 56.66 37.51 ;
      RECT  55.77 37.51 58.85 37.81 ;
      RECT  56.15 42.25 56.63 42.16 ;
      RECT  55.77 42.16 58.85 41.86 ;
      RECT  56.15 41.86 56.64 41.76 ;
      RECT  56.13 38.04 56.66 37.81 ;
      RECT  55.77 37.81 58.85 37.51 ;
      RECT  56.15 41.77 56.63 41.86 ;
      RECT  55.77 41.86 58.85 42.16 ;
      RECT  56.15 42.16 56.64 42.26 ;
      RECT  56.13 45.98 56.66 46.21 ;
      RECT  55.77 46.21 58.85 46.51 ;
      RECT  56.15 50.95 56.63 50.86 ;
      RECT  55.77 50.86 58.85 50.56 ;
      RECT  56.15 50.56 56.64 50.46 ;
      RECT  56.13 46.74 56.66 46.51 ;
      RECT  55.77 46.51 58.85 46.21 ;
      RECT  56.15 50.47 56.63 50.56 ;
      RECT  55.77 50.56 58.85 50.86 ;
      RECT  56.15 50.86 56.64 50.96 ;
      RECT  56.13 54.68 56.66 54.91 ;
      RECT  55.77 54.91 58.85 55.21 ;
      RECT  56.15 59.65 56.63 59.56 ;
      RECT  55.77 59.56 58.85 59.26 ;
      RECT  56.15 59.26 56.64 59.16 ;
      RECT  56.13 55.44 56.66 55.21 ;
      RECT  55.77 55.21 58.85 54.91 ;
      RECT  56.15 59.17 56.63 59.26 ;
      RECT  55.77 59.26 58.85 59.56 ;
      RECT  56.15 59.56 56.64 59.66 ;
      RECT  56.13 63.38 56.66 63.61 ;
      RECT  55.77 63.61 58.85 63.91 ;
      RECT  56.15 68.35 56.63 68.26 ;
      RECT  55.77 68.26 58.85 67.96 ;
      RECT  56.15 67.96 56.64 67.86 ;
      RECT  56.13 64.14 56.66 63.91 ;
      RECT  55.77 63.91 58.85 63.61 ;
      RECT  56.15 67.87 56.63 67.96 ;
      RECT  55.77 67.96 58.85 68.26 ;
      RECT  56.15 68.26 56.64 68.36 ;
      RECT  56.13 72.08 56.66 72.31 ;
      RECT  55.77 72.31 58.85 72.61 ;
      RECT  56.15 77.05 56.63 76.96 ;
      RECT  55.77 76.96 58.85 76.66 ;
      RECT  56.15 76.66 56.64 76.56 ;
      RECT  56.13 72.84 56.66 72.61 ;
      RECT  55.77 72.61 58.85 72.31 ;
      RECT  56.15 76.57 56.63 76.66 ;
      RECT  55.77 76.66 58.85 76.96 ;
      RECT  56.15 76.96 56.64 77.06 ;
      RECT  56.13 80.78 56.66 81.01 ;
      RECT  55.77 81.01 58.85 81.31 ;
      RECT  56.15 85.75 56.63 85.66 ;
      RECT  55.77 85.66 58.85 85.36 ;
      RECT  56.15 85.36 56.64 85.26 ;
      RECT  56.13 81.54 56.66 81.31 ;
      RECT  55.77 81.31 58.85 81.01 ;
      RECT  56.15 85.27 56.63 85.36 ;
      RECT  55.77 85.36 58.85 85.66 ;
      RECT  56.15 85.66 56.64 85.76 ;
      RECT  56.13 89.48 56.66 89.71 ;
      RECT  55.77 89.71 58.85 90.01 ;
      RECT  56.15 94.45 56.63 94.36 ;
      RECT  55.77 94.36 58.85 94.06 ;
      RECT  56.15 94.06 56.64 93.96 ;
      RECT  56.13 90.24 56.66 90.01 ;
      RECT  55.77 90.01 58.85 89.71 ;
      RECT  56.15 93.97 56.63 94.06 ;
      RECT  55.77 94.06 58.85 94.36 ;
      RECT  56.15 94.36 56.64 94.46 ;
      RECT  56.13 98.18 56.66 98.41 ;
      RECT  55.77 98.41 58.85 98.71 ;
      RECT  56.15 103.15 56.63 103.06 ;
      RECT  55.77 103.06 58.85 102.76 ;
      RECT  56.15 102.76 56.64 102.66 ;
      RECT  56.13 98.94 56.66 98.71 ;
      RECT  55.77 98.71 58.85 98.41 ;
      RECT  56.15 102.67 56.63 102.76 ;
      RECT  55.77 102.76 58.85 103.06 ;
      RECT  56.15 103.06 56.64 103.16 ;
      RECT  56.13 106.88 56.66 107.11 ;
      RECT  55.77 107.11 58.85 107.41 ;
      RECT  55.77 98.41 58.85 98.71 ;
      RECT  55.77 98.41 58.85 98.71 ;
      RECT  55.77 54.91 58.85 55.21 ;
      RECT  55.77 46.21 58.85 46.51 ;
      RECT  55.77 63.61 58.85 63.91 ;
      RECT  55.77 37.51 58.85 37.81 ;
      RECT  55.77 37.51 58.85 37.81 ;
      RECT  55.77 28.81 58.85 29.11 ;
      RECT  55.77 28.81 58.85 29.11 ;
      RECT  55.77 72.31 58.85 72.61 ;
      RECT  55.77 81.01 58.85 81.31 ;
      RECT  55.77 81.01 58.85 81.31 ;
      RECT  55.77 107.11 58.85 107.41 ;
      RECT  55.77 89.71 58.85 90.01 ;
      RECT  55.77 63.61 58.85 63.91 ;
      RECT  55.77 89.71 58.85 90.01 ;
      RECT  55.77 54.91 58.85 55.21 ;
      RECT  55.77 85.36 58.85 85.66 ;
      RECT  55.77 41.86 58.85 42.16 ;
      RECT  55.77 33.16 58.85 33.46 ;
      RECT  55.77 50.56 58.85 50.86 ;
      RECT  55.77 76.66 58.85 76.96 ;
      RECT  55.77 24.46 58.85 24.76 ;
      RECT  55.77 94.06 58.85 94.36 ;
      RECT  55.77 59.26 58.85 59.56 ;
      RECT  55.77 102.76 58.85 103.06 ;
      RECT  55.77 67.96 58.85 68.26 ;
      RECT  44.84 54.91 45.14 55.21 ;
      RECT  46.53 81.01 49.61 81.31 ;
      RECT  57.16 63.61 57.46 63.91 ;
      RECT  47.92 28.81 48.22 29.11 ;
      RECT  46.53 46.21 49.61 46.51 ;
      RECT  57.16 54.91 57.46 55.21 ;
      RECT  44.84 46.21 45.14 46.51 ;
      RECT  57.16 46.21 57.46 46.51 ;
      RECT  46.53 98.41 49.61 98.71 ;
      RECT  46.53 89.71 49.61 90.01 ;
      RECT  44.84 89.71 45.14 90.01 ;
      RECT  57.16 72.31 57.46 72.61 ;
      RECT  51.0 28.81 51.3 29.11 ;
      RECT  54.08 107.11 54.38 107.41 ;
      RECT  57.16 37.51 57.46 37.81 ;
      RECT  57.16 89.71 57.46 90.01 ;
      RECT  46.53 54.91 49.61 55.21 ;
      RECT  46.53 63.61 49.61 63.91 ;
      RECT  44.84 81.01 45.14 81.31 ;
      RECT  54.08 28.81 54.38 29.11 ;
      RECT  57.16 28.81 57.46 29.11 ;
      RECT  44.84 63.61 45.14 63.91 ;
      RECT  46.53 37.51 49.61 37.81 ;
      RECT  57.16 98.41 57.46 98.71 ;
      RECT  44.84 28.81 45.14 29.11 ;
      RECT  57.16 107.11 57.46 107.41 ;
      RECT  44.84 72.31 45.14 72.61 ;
      RECT  51.0 107.11 51.3 107.41 ;
      RECT  57.16 81.01 57.46 81.31 ;
      RECT  47.92 107.11 48.22 107.41 ;
      RECT  44.84 98.41 45.14 98.71 ;
      RECT  44.84 107.11 45.14 107.41 ;
      RECT  46.53 72.31 49.61 72.61 ;
      RECT  46.53 28.81 49.61 29.11 ;
      RECT  44.84 37.51 45.14 37.81 ;
      RECT  44.84 67.96 45.14 68.26 ;
      RECT  47.92 102.76 48.22 103.06 ;
      RECT  46.53 102.76 49.61 103.06 ;
      RECT  44.84 85.36 45.14 85.66 ;
      RECT  46.53 33.16 49.61 33.46 ;
      RECT  44.84 102.76 45.14 103.06 ;
      RECT  57.16 41.86 57.46 42.16 ;
      RECT  57.16 76.66 57.46 76.96 ;
      RECT  44.84 94.06 45.14 94.36 ;
      RECT  54.08 102.76 54.38 103.06 ;
      RECT  46.53 59.26 49.61 59.56 ;
      RECT  44.84 76.66 45.14 76.96 ;
      RECT  46.53 76.66 49.61 76.96 ;
      RECT  42.29 24.755 42.81 25.275 ;
      RECT  42.29 103.055 42.81 103.575 ;
      RECT  59.49 24.755 60.01 25.275 ;
      RECT  51.0 24.46 51.3 24.76 ;
      RECT  44.84 24.46 45.14 24.76 ;
      RECT  57.16 85.36 57.46 85.66 ;
      RECT  57.16 67.96 57.46 68.26 ;
      RECT  57.16 102.76 57.46 103.06 ;
      RECT  47.92 24.46 48.22 24.76 ;
      RECT  44.84 59.26 45.14 59.56 ;
      RECT  57.16 33.16 57.46 33.46 ;
      RECT  54.08 24.46 54.38 24.76 ;
      RECT  59.49 103.055 60.01 103.575 ;
      RECT  57.16 50.56 57.46 50.86 ;
      RECT  46.53 41.86 49.61 42.16 ;
      RECT  51.0 102.76 51.3 103.06 ;
      RECT  46.53 67.96 49.61 68.26 ;
      RECT  46.53 94.06 49.61 94.36 ;
      RECT  44.84 50.56 45.14 50.86 ;
      RECT  46.53 85.36 49.61 85.66 ;
      RECT  57.16 59.26 57.46 59.56 ;
      RECT  57.16 24.46 57.46 24.76 ;
      RECT  46.53 50.56 49.61 50.86 ;
      RECT  57.16 94.06 57.46 94.36 ;
      RECT  44.84 41.86 45.14 42.16 ;
      RECT  44.84 33.16 45.14 33.46 ;
      RECT  48.365 21.9 48.885 22.42 ;
      RECT  51.445 21.9 51.965 22.42 ;
      RECT  54.525 21.9 55.045 22.42 ;
      RECT  51.445 21.9 51.965 22.42 ;
      RECT  54.525 21.9 55.045 22.42 ;
      RECT  48.365 21.9 48.885 22.42 ;
      RECT  49.61 13.47 52.69 13.82 ;
      RECT  49.61 8.91 52.69 9.21 ;
      RECT  49.8 13.38 50.33 13.47 ;
      RECT  49.91 8.81 50.43 8.91 ;
      RECT  49.8 13.82 50.33 13.91 ;
      RECT  49.91 9.21 50.43 9.31 ;
      RECT  52.69 13.47 55.77 13.82 ;
      RECT  52.69 8.91 55.77 9.21 ;
      RECT  52.88 13.38 53.41 13.47 ;
      RECT  52.99 8.81 53.51 8.91 ;
      RECT  52.88 13.82 53.41 13.91 ;
      RECT  52.99 9.21 53.51 9.31 ;
      RECT  54.08 13.495 54.38 13.795 ;
      RECT  51.0 13.495 51.3 13.795 ;
      RECT  51.0 8.91 51.3 9.21 ;
      RECT  54.08 8.91 54.38 9.21 ;
      RECT  49.61 -0.17 52.69 0.18 ;
      RECT  51.47 4.46 51.92 4.51 ;
      RECT  51.47 4.06 51.92 4.11 ;
      RECT  51.29 6.84 51.78 6.9 ;
      RECT  51.36 0.18 51.87 0.26 ;
      RECT  49.61 4.11 52.69 4.46 ;
      RECT  49.61 6.9 52.69 7.25 ;
      RECT  51.29 7.25 51.78 7.33 ;
      RECT  51.36 -0.25 51.87 -0.17 ;
      RECT  52.69 -0.17 55.77 0.18 ;
      RECT  54.55 4.46 55.0 4.51 ;
      RECT  54.55 4.06 55.0 4.11 ;
      RECT  54.37 6.84 54.86 6.9 ;
      RECT  54.44 0.18 54.95 0.26 ;
      RECT  52.69 4.11 55.77 4.46 ;
      RECT  52.69 6.9 55.77 7.25 ;
      RECT  54.37 7.25 54.86 7.33 ;
      RECT  54.44 -0.25 54.95 -0.17 ;
      RECT  54.08 4.135 54.38 4.435 ;
      RECT  51.0 4.135 51.3 4.435 ;
      RECT  51.0 6.925 51.3 7.225 ;
      RECT  54.08 6.925 54.38 7.225 ;
      RECT  51.0 -0.145 51.3 0.155 ;
      RECT  54.08 -0.145 54.38 0.155 ;
      RECT  54.08 4.435 54.38 4.135 ;
      RECT  54.525 22.42 55.045 21.9 ;
      RECT  51.0 13.795 51.3 13.495 ;
      RECT  51.0 4.435 51.3 4.135 ;
      RECT  48.365 22.42 48.885 21.9 ;
      RECT  51.445 22.42 51.965 21.9 ;
      RECT  54.08 13.795 54.38 13.495 ;
      RECT  54.08 9.21 54.38 8.91 ;
      RECT  51.0 0.155 51.3 -0.145 ;
      RECT  51.0 9.21 51.3 8.91 ;
      RECT  54.08 7.225 54.38 6.925 ;
      RECT  54.08 0.155 54.38 -0.145 ;
      RECT  51.0 7.225 51.3 6.925 ;
      RECT  5.18 37.4 5.7 37.92 ;
      RECT  5.18 37.4 5.7 37.92 ;
      RECT  12.28 46.1 12.8 46.62 ;
      RECT  5.18 46.1 5.7 46.62 ;
      RECT  12.28 37.4 12.8 37.92 ;
      RECT  12.28 37.4 12.8 37.92 ;
      RECT  12.28 50.45 12.8 50.97 ;
      RECT  5.18 50.45 5.7 50.97 ;
      RECT  12.28 41.75 12.8 42.27 ;
      RECT  12.28 33.05 12.8 33.57 ;
      RECT  5.18 41.75 5.7 42.27 ;
      RECT  5.18 33.05 5.7 33.57 ;
      RECT  5.18 63.5 5.7 64.02 ;
      RECT  5.18 63.5 5.7 64.02 ;
      RECT  12.28 72.2 12.8 72.72 ;
      RECT  5.18 72.2 5.7 72.72 ;
      RECT  12.28 63.5 12.8 64.02 ;
      RECT  12.28 63.5 12.8 64.02 ;
      RECT  12.28 76.55 12.8 77.07 ;
      RECT  5.18 76.55 5.7 77.07 ;
      RECT  12.28 67.85 12.8 68.37 ;
      RECT  12.28 59.15 12.8 59.67 ;
      RECT  5.18 67.85 5.7 68.37 ;
      RECT  5.18 59.15 5.7 59.67 ;
      RECT  12.28 63.5 12.8 64.02 ;
      RECT  12.28 37.4 12.8 37.92 ;
      RECT  32.17 89.6 32.69 90.12 ;
      RECT  32.17 89.6 32.69 90.12 ;
      RECT  32.17 72.2 32.69 72.72 ;
      RECT  32.17 72.2 32.69 72.72 ;
      RECT  32.17 80.9 32.69 81.42 ;
      RECT  5.18 72.2 5.7 72.72 ;
      RECT  32.17 37.4 32.69 37.92 ;
      RECT  5.18 46.1 5.7 46.62 ;
      RECT  32.17 54.8 32.69 55.32 ;
      RECT  5.18 63.5 5.7 64.02 ;
      RECT  12.28 46.1 12.8 46.62 ;
      RECT  32.17 46.1 32.69 46.62 ;
      RECT  32.17 98.3 32.69 98.82 ;
      RECT  12.28 72.2 12.8 72.72 ;
      RECT  5.18 37.4 5.7 37.92 ;
      RECT  32.17 63.5 32.69 64.02 ;
      RECT  32.17 37.4 32.69 37.92 ;
      RECT  32.17 93.95 32.69 94.47 ;
      RECT  12.28 50.45 12.8 50.97 ;
      RECT  32.17 76.55 32.69 77.07 ;
      RECT  12.28 67.85 12.8 68.37 ;
      RECT  32.17 59.15 32.69 59.67 ;
      RECT  32.17 102.65 32.69 103.17 ;
      RECT  32.17 67.85 32.69 68.37 ;
      RECT  5.18 59.15 5.7 59.67 ;
      RECT  12.28 59.15 12.8 59.67 ;
      RECT  32.17 85.25 32.69 85.77 ;
      RECT  12.28 33.05 12.8 33.57 ;
      RECT  32.17 41.75 32.69 42.27 ;
      RECT  5.18 50.45 5.7 50.97 ;
      RECT  12.28 41.75 12.8 42.27 ;
      RECT  5.18 76.55 5.7 77.07 ;
      RECT  12.28 76.55 12.8 77.07 ;
      RECT  32.17 50.45 32.69 50.97 ;
      RECT  32.17 33.05 32.69 33.57 ;
      RECT  5.18 41.75 5.7 42.27 ;
      RECT  5.18 33.05 5.7 33.57 ;
      RECT  5.18 67.85 5.7 68.37 ;
      RECT  39.04 72.2 39.56 72.72 ;
      RECT  39.04 54.8 39.56 55.32 ;
      RECT  39.04 72.2 39.56 72.72 ;
      RECT  39.04 46.1 39.56 46.62 ;
      RECT  39.04 98.3 39.56 98.82 ;
      RECT  39.04 37.4 39.56 37.92 ;
      RECT  39.04 37.4 39.56 37.92 ;
      RECT  39.04 63.5 39.56 64.02 ;
      RECT  39.04 89.6 39.56 90.12 ;
      RECT  39.04 89.6 39.56 90.12 ;
      RECT  39.04 80.9 39.56 81.42 ;
      RECT  39.04 93.95 39.56 94.47 ;
      RECT  39.04 76.55 39.56 77.07 ;
      RECT  39.04 59.15 39.56 59.67 ;
      RECT  39.04 102.65 39.56 103.17 ;
      RECT  39.04 50.45 39.56 50.97 ;
      RECT  39.04 85.25 39.56 85.77 ;
      RECT  39.04 41.75 39.56 42.27 ;
      RECT  39.04 67.85 39.56 68.37 ;
      RECT  39.04 33.05 39.56 33.57 ;
      RECT  39.04 80.9 39.56 81.42 ;
      RECT  32.17 63.5 32.69 64.02 ;
      RECT  39.04 89.6 39.56 90.12 ;
      RECT  5.18 37.4 5.7 37.92 ;
      RECT  12.28 72.2 12.8 72.72 ;
      RECT  39.04 98.3 39.56 98.82 ;
      RECT  5.18 63.5 5.7 64.02 ;
      RECT  5.18 46.1 5.7 46.62 ;
      RECT  32.17 37.4 32.69 37.92 ;
      RECT  32.17 98.3 32.69 98.82 ;
      RECT  39.04 72.2 39.56 72.72 ;
      RECT  32.17 46.1 32.69 46.62 ;
      RECT  12.28 63.5 12.8 64.02 ;
      RECT  32.17 80.9 32.69 81.42 ;
      RECT  39.04 63.5 39.56 64.02 ;
      RECT  39.04 54.8 39.56 55.32 ;
      RECT  32.69 29.895 33.21 30.415 ;
      RECT  5.18 72.2 5.7 72.72 ;
      RECT  32.17 72.2 32.69 72.72 ;
      RECT  32.17 89.6 32.69 90.12 ;
      RECT  32.17 54.8 32.69 55.32 ;
      RECT  32.17 28.7 32.69 29.22 ;
      RECT  39.04 46.1 39.56 46.62 ;
      RECT  12.28 37.4 12.8 37.92 ;
      RECT  39.04 37.4 39.56 37.92 ;
      RECT  12.28 46.1 12.8 46.62 ;
      RECT  32.17 59.15 32.69 59.67 ;
      RECT  32.17 93.95 32.69 94.47 ;
      RECT  5.18 41.75 5.7 42.27 ;
      RECT  39.04 76.55 39.56 77.07 ;
      RECT  32.17 33.05 32.69 33.57 ;
      RECT  5.18 76.55 5.7 77.07 ;
      RECT  39.04 93.95 39.56 94.47 ;
      RECT  12.28 50.45 12.8 50.97 ;
      RECT  39.04 33.05 39.56 33.57 ;
      RECT  5.18 59.15 5.7 59.67 ;
      RECT  32.17 67.85 32.69 68.37 ;
      RECT  39.04 102.65 39.56 103.17 ;
      RECT  32.17 102.65 32.69 103.17 ;
      RECT  12.28 33.05 12.8 33.57 ;
      RECT  12.28 59.15 12.8 59.67 ;
      RECT  39.04 67.85 39.56 68.37 ;
      RECT  12.28 76.55 12.8 77.07 ;
      RECT  32.17 76.55 32.69 77.07 ;
      RECT  39.04 85.25 39.56 85.77 ;
      RECT  12.28 41.75 12.8 42.27 ;
      RECT  39.04 41.75 39.56 42.27 ;
      RECT  32.17 41.75 32.69 42.27 ;
      RECT  32.17 85.25 32.69 85.77 ;
      RECT  12.28 67.85 12.8 68.37 ;
      RECT  32.17 50.45 32.69 50.97 ;
      RECT  5.18 50.45 5.7 50.97 ;
      RECT  5.18 67.85 5.7 68.37 ;
      RECT  39.04 59.15 39.56 59.67 ;
      RECT  5.18 33.05 5.7 33.57 ;
      RECT  39.04 50.45 39.56 50.97 ;
      RECT  0.0 14.66 47.19 14.96 ;
      RECT  54.08 13.495 54.38 13.795 ;
      RECT  44.84 54.91 45.14 55.21 ;
      RECT  46.53 81.01 49.61 81.31 ;
      RECT  57.16 63.61 57.46 63.91 ;
      RECT  5.18 63.5 5.7 64.02 ;
      RECT  47.92 28.81 48.22 29.11 ;
      RECT  32.17 89.6 32.69 90.12 ;
      RECT  46.53 46.21 49.61 46.51 ;
      RECT  12.28 37.4 12.8 37.92 ;
      RECT  57.16 54.91 57.46 55.21 ;
      RECT  44.84 46.21 45.14 46.51 ;
      RECT  5.18 46.1 5.7 46.62 ;
      RECT  57.16 46.21 57.46 46.51 ;
      RECT  12.28 63.5 12.8 64.02 ;
      RECT  39.04 80.9 39.56 81.42 ;
      RECT  46.53 98.41 49.61 98.71 ;
      RECT  46.53 89.71 49.61 90.01 ;
      RECT  51.0 13.495 51.3 13.795 ;
      RECT  44.84 89.71 45.14 90.01 ;
      RECT  12.28 46.1 12.8 46.62 ;
      RECT  51.445 21.9 51.965 22.42 ;
      RECT  32.17 80.9 32.69 81.42 ;
      RECT  57.16 72.31 57.46 72.61 ;
      RECT  51.0 28.81 51.3 29.11 ;
      RECT  32.17 37.4 32.69 37.92 ;
      RECT  32.17 46.1 32.69 46.62 ;
      RECT  32.69 29.895 33.21 30.415 ;
      RECT  5.18 72.2 5.7 72.72 ;
      RECT  39.04 46.1 39.56 46.62 ;
      RECT  54.08 107.11 54.38 107.41 ;
      RECT  57.16 89.71 57.46 90.01 ;
      RECT  46.53 54.91 49.61 55.21 ;
      RECT  57.16 37.51 57.46 37.81 ;
      RECT  46.53 63.61 49.61 63.91 ;
      RECT  44.84 81.01 45.14 81.31 ;
      RECT  51.0 4.135 51.3 4.435 ;
      RECT  32.17 54.8 32.69 55.32 ;
      RECT  39.04 63.5 39.56 64.02 ;
      RECT  54.08 28.81 54.38 29.11 ;
      RECT  32.17 63.5 32.69 64.02 ;
      RECT  57.16 28.81 57.46 29.11 ;
      RECT  44.84 63.61 45.14 63.91 ;
      RECT  46.53 37.51 49.61 37.81 ;
      RECT  57.16 98.41 57.46 98.71 ;
      RECT  44.84 28.81 45.14 29.11 ;
      RECT  57.16 107.11 57.46 107.41 ;
      RECT  39.04 54.8 39.56 55.32 ;
      RECT  48.365 21.9 48.885 22.42 ;
      RECT  44.84 72.31 45.14 72.61 ;
      RECT  51.0 107.11 51.3 107.41 ;
      RECT  57.16 81.01 57.46 81.31 ;
      RECT  39.04 37.4 39.56 37.92 ;
      RECT  32.17 72.2 32.69 72.72 ;
      RECT  47.92 107.11 48.22 107.41 ;
      RECT  54.525 21.9 55.045 22.42 ;
      RECT  44.84 98.41 45.14 98.71 ;
      RECT  5.18 37.4 5.7 37.92 ;
      RECT  32.17 28.7 32.69 29.22 ;
      RECT  39.04 89.6 39.56 90.12 ;
      RECT  39.04 98.3 39.56 98.82 ;
      RECT  32.17 98.3 32.69 98.82 ;
      RECT  44.84 107.11 45.14 107.41 ;
      RECT  39.04 72.2 39.56 72.72 ;
      RECT  46.53 72.31 49.61 72.61 ;
      RECT  46.53 28.81 49.61 29.11 ;
      RECT  44.84 37.51 45.14 37.81 ;
      RECT  12.28 72.2 12.8 72.72 ;
      RECT  54.08 4.135 54.38 4.435 ;
      RECT  44.84 67.96 45.14 68.26 ;
      RECT  47.92 102.76 48.22 103.06 ;
      RECT  46.53 102.76 49.61 103.06 ;
      RECT  39.04 41.75 39.56 42.27 ;
      RECT  46.53 33.16 49.61 33.46 ;
      RECT  44.84 85.36 45.14 85.66 ;
      RECT  39.04 59.15 39.56 59.67 ;
      RECT  39.04 50.45 39.56 50.97 ;
      RECT  44.84 102.76 45.14 103.06 ;
      RECT  57.16 41.86 57.46 42.16 ;
      RECT  57.16 76.66 57.46 76.96 ;
      RECT  44.84 94.06 45.14 94.36 ;
      RECT  54.08 102.76 54.38 103.06 ;
      RECT  32.17 85.25 32.69 85.77 ;
      RECT  32.17 93.95 32.69 94.47 ;
      RECT  46.53 59.26 49.61 59.56 ;
      RECT  12.28 41.75 12.8 42.27 ;
      RECT  39.04 33.05 39.56 33.57 ;
      RECT  39.04 67.85 39.56 68.37 ;
      RECT  5.18 33.05 5.7 33.57 ;
      RECT  44.84 76.66 45.14 76.96 ;
      RECT  46.53 76.66 49.61 76.96 ;
      RECT  12.28 50.45 12.8 50.97 ;
      RECT  42.29 24.755 42.81 25.275 ;
      RECT  51.0 8.91 51.3 9.21 ;
      RECT  42.29 103.055 42.81 103.575 ;
      RECT  59.49 24.755 60.01 25.275 ;
      RECT  54.08 8.91 54.38 9.21 ;
      RECT  51.0 24.46 51.3 24.76 ;
      RECT  32.17 102.65 32.69 103.17 ;
      RECT  32.17 67.85 32.69 68.37 ;
      RECT  44.84 24.46 45.14 24.76 ;
      RECT  32.17 50.45 32.69 50.97 ;
      RECT  57.16 85.36 57.46 85.66 ;
      RECT  32.17 76.55 32.69 77.07 ;
      RECT  57.16 67.96 57.46 68.26 ;
      RECT  57.16 102.76 57.46 103.06 ;
      RECT  47.92 24.46 48.22 24.76 ;
      RECT  44.84 59.26 45.14 59.56 ;
      RECT  5.18 41.75 5.7 42.27 ;
      RECT  5.18 59.15 5.7 59.67 ;
      RECT  39.04 76.55 39.56 77.07 ;
      RECT  39.04 102.65 39.56 103.17 ;
      RECT  32.17 41.75 32.69 42.27 ;
      RECT  57.16 33.16 57.46 33.46 ;
      RECT  32.17 33.05 32.69 33.57 ;
      RECT  12.28 33.05 12.8 33.57 ;
      RECT  12.28 59.15 12.8 59.67 ;
      RECT  54.08 24.46 54.38 24.76 ;
      RECT  59.49 103.055 60.01 103.575 ;
      RECT  5.18 50.45 5.7 50.97 ;
      RECT  57.16 50.56 57.46 50.86 ;
      RECT  54.08 6.925 54.38 7.225 ;
      RECT  46.53 41.86 49.61 42.16 ;
      RECT  5.18 67.85 5.7 68.37 ;
      RECT  51.0 102.76 51.3 103.06 ;
      RECT  39.04 93.95 39.56 94.47 ;
      RECT  46.53 67.96 49.61 68.26 ;
      RECT  51.0 -0.145 51.3 0.155 ;
      RECT  54.08 -0.145 54.38 0.155 ;
      RECT  46.53 94.06 49.61 94.36 ;
      RECT  44.84 50.56 45.14 50.86 ;
      RECT  46.53 85.36 49.61 85.66 ;
      RECT  12.28 76.55 12.8 77.07 ;
      RECT  57.16 59.26 57.46 59.56 ;
      RECT  57.16 24.46 57.46 24.76 ;
      RECT  46.53 50.56 49.61 50.86 ;
      RECT  51.0 6.925 51.3 7.225 ;
      RECT  32.17 59.15 32.69 59.67 ;
      RECT  12.28 67.85 12.8 68.37 ;
      RECT  57.16 94.06 57.46 94.36 ;
      RECT  44.84 41.86 45.14 42.16 ;
      RECT  39.04 85.25 39.56 85.77 ;
      RECT  5.18 76.55 5.7 77.07 ;
      RECT  44.84 33.16 45.14 33.46 ;
      RECT  -55.65 -5.475 -55.13 -4.955 ;
      RECT  -55.65 -5.485 -55.13 -4.965 ;
      RECT  -55.71 -1.385 -55.19 -0.865 ;
      RECT  -55.71 -9.575 -55.19 -9.055 ;
      RECT  -45.17 32.75 -45.69 33.27 ;
      RECT  -45.17 32.75 -45.69 33.27 ;
      RECT  -51.45 66.35 -51.97 66.87 ;
      RECT  -51.45 83.15 -51.97 83.67 ;
      RECT  -51.45 99.95 -51.97 100.47 ;
      RECT  -45.17 83.15 -45.69 83.67 ;
      RECT  -45.17 83.15 -45.69 83.67 ;
      RECT  -51.45 32.75 -51.97 33.27 ;
      RECT  -51.45 32.75 -51.97 33.27 ;
      RECT  -51.45 49.55 -51.97 50.07 ;
      RECT  -45.17 66.35 -45.69 66.87 ;
      RECT  -45.17 99.95 -45.69 100.47 ;
      RECT  -51.45 83.15 -51.97 83.67 ;
      RECT  -45.17 49.55 -45.69 50.07 ;
      RECT  -45.17 57.95 -45.69 58.47 ;
      RECT  -51.45 41.15 -51.97 41.67 ;
      RECT  -51.45 57.95 -51.97 58.47 ;
      RECT  -45.17 91.55 -45.69 92.07 ;
      RECT  -45.17 74.75 -45.69 75.27 ;
      RECT  -51.45 74.75 -51.97 75.27 ;
      RECT  -51.45 24.35 -51.97 24.87 ;
      RECT  -45.17 41.15 -45.69 41.67 ;
      RECT  -51.45 91.55 -51.97 92.07 ;
      RECT  -45.17 24.35 -45.69 24.87 ;
      RECT  -45.69 66.35 -45.17 66.87 ;
      RECT  -51.97 49.55 -51.45 50.07 ;
      RECT  -45.69 99.95 -45.17 100.47 ;
      RECT  -45.69 49.55 -45.17 50.07 ;
      RECT  -45.69 32.75 -45.17 33.27 ;
      RECT  -51.97 83.15 -51.45 83.67 ;
      RECT  -55.65 -5.475 -55.13 -4.955 ;
      RECT  -51.97 32.75 -51.45 33.27 ;
      RECT  -51.97 66.35 -51.45 66.87 ;
      RECT  -45.69 83.15 -45.17 83.67 ;
      RECT  -51.97 99.95 -51.45 100.47 ;
      RECT  -55.65 -5.485 -55.13 -4.965 ;
      RECT  -51.97 91.55 -51.45 92.07 ;
      RECT  -51.97 24.35 -51.45 24.87 ;
      RECT  -45.69 57.95 -45.17 58.47 ;
      RECT  -51.97 74.75 -51.45 75.27 ;
      RECT  -55.71 -1.385 -55.19 -0.865 ;
      RECT  -45.69 91.55 -45.17 92.07 ;
      RECT  -45.69 74.75 -45.17 75.27 ;
      RECT  -51.97 57.95 -51.45 58.47 ;
      RECT  -45.69 41.15 -45.17 41.67 ;
      RECT  -45.69 24.35 -45.17 24.87 ;
      RECT  -51.97 41.15 -51.45 41.67 ;
      RECT  -55.71 -9.575 -55.19 -9.055 ;
      RECT  -14.03 103.2 -1.32 103.5 ;
      RECT  -7.905 113.425 -7.385 113.945 ;
      RECT  -7.905 105.245 -7.385 105.765 ;
      RECT  -7.905 113.415 -7.385 113.935 ;
      RECT  -7.905 105.235 -7.385 105.755 ;
      RECT  -8.025 109.325 -7.505 109.845 ;
      RECT  -8.025 101.145 -7.505 101.665 ;
      RECT  -8.025 117.515 -7.505 118.035 ;
      RECT  -8.025 109.335 -7.505 109.855 ;
      RECT  11.39 -7.52 36.81 -7.22 ;
      RECT  17.515 -5.485 18.035 -4.965 ;
      RECT  30.225 -5.485 30.745 -4.965 ;
      RECT  17.395 -9.575 17.915 -9.055 ;
      RECT  30.105 -9.575 30.625 -9.055 ;
   LAYER  m4 ;
   END
   END    sram_2_16_sky130A
END    LIBRARY
