magic
tech sky130A
timestamp 1616584750
<< nwell >>
rect 0 376 260 558
<< nmos >>
rect 53 153 68 279
rect 195 153 210 279
rect 76 104 118 119
rect 145 104 187 119
<< pmos >>
rect 53 404 68 459
rect 186 404 201 459
<< ndiff >>
rect 18 271 53 279
rect 18 254 26 271
rect 43 254 53 271
rect 18 226 53 254
rect 18 209 26 226
rect 43 209 53 226
rect 18 178 53 209
rect 18 161 26 178
rect 43 161 53 178
rect 18 153 53 161
rect 68 271 118 279
rect 68 254 93 271
rect 110 254 118 271
rect 68 178 118 254
rect 68 161 93 178
rect 110 161 118 178
rect 68 153 118 161
rect 76 119 118 153
rect 145 271 195 279
rect 145 254 153 271
rect 170 254 195 271
rect 145 178 195 254
rect 145 161 153 178
rect 170 161 195 178
rect 145 153 195 161
rect 210 271 245 279
rect 210 254 220 271
rect 237 254 245 271
rect 210 229 245 254
rect 210 212 220 229
rect 237 212 245 229
rect 210 178 245 212
rect 210 161 220 178
rect 237 161 245 178
rect 210 153 245 161
rect 145 119 187 153
rect 76 94 118 104
rect 76 77 93 94
rect 110 77 118 94
rect 76 70 118 77
rect 145 95 187 104
rect 145 78 153 95
rect 170 78 187 95
rect 145 70 187 78
<< pdiff >>
rect 18 451 53 459
rect 18 434 26 451
rect 43 434 53 451
rect 18 404 53 434
rect 68 429 103 459
rect 68 412 78 429
rect 95 412 103 429
rect 68 404 103 412
rect 151 451 186 459
rect 151 434 159 451
rect 176 434 186 451
rect 151 404 186 434
rect 201 429 236 459
rect 201 412 211 429
rect 228 412 236 429
rect 201 404 236 412
<< ndiffc >>
rect 26 254 43 271
rect 26 209 43 226
rect 26 161 43 178
rect 93 254 110 271
rect 93 161 110 178
rect 153 254 170 271
rect 153 161 170 178
rect 220 254 237 271
rect 220 212 237 229
rect 220 161 237 178
rect 93 77 110 94
rect 153 78 170 95
<< pdiffc >>
rect 26 434 43 451
rect 78 412 95 429
rect 159 434 176 451
rect 211 412 228 429
<< psubdiff >>
rect 7 9 48 21
rect 7 -8 19 9
rect 36 -8 48 9
rect 7 -20 48 -8
<< nsubdiff >>
rect 18 521 71 539
rect 18 504 36 521
rect 53 504 71 521
rect 18 486 71 504
<< psubdiffcont >>
rect 19 -8 36 9
<< nsubdiffcont >>
rect 36 504 53 521
<< poly >>
rect 53 459 68 472
rect 186 459 201 472
rect 53 383 68 404
rect 53 375 165 383
rect 53 368 140 375
rect 53 279 68 368
rect 132 358 140 368
rect 157 358 165 375
rect 132 350 165 358
rect 90 321 123 329
rect 90 304 98 321
rect 115 318 123 321
rect 186 318 201 404
rect 115 304 210 318
rect 90 303 210 304
rect 90 296 123 303
rect 195 279 210 303
rect 53 140 68 153
rect 195 140 210 153
rect 0 111 76 119
rect 0 104 26 111
rect 18 94 26 104
rect 43 104 76 111
rect 118 104 145 119
rect 187 104 260 119
rect 43 94 51 104
rect 18 86 51 94
<< polycont >>
rect 140 358 157 375
rect 98 304 115 321
rect 26 94 43 111
<< locali >>
rect 28 521 61 529
rect 0 504 36 521
rect 53 504 127 521
rect 144 504 260 521
rect 28 496 61 504
rect 28 459 45 496
rect 18 451 51 459
rect 18 434 26 451
rect 43 434 51 451
rect 151 451 184 459
rect 18 426 51 434
rect 70 429 103 437
rect 70 412 78 429
rect 95 412 103 429
rect 70 404 103 412
rect 151 434 159 451
rect 176 434 184 451
rect 211 437 228 504
rect 151 426 184 434
rect 203 429 236 437
rect 85 329 102 404
rect 151 383 168 426
rect 203 412 211 429
rect 228 412 236 429
rect 203 404 236 412
rect 132 375 168 383
rect 132 358 140 375
rect 157 358 168 375
rect 132 350 168 358
rect 85 321 123 329
rect 85 304 98 321
rect 115 304 123 321
rect 85 296 123 304
rect 85 279 102 296
rect 151 279 168 350
rect 18 271 51 279
rect 18 254 26 271
rect 43 254 51 271
rect 18 226 51 254
rect 85 271 118 279
rect 85 254 93 271
rect 110 254 118 271
rect 85 246 118 254
rect 145 271 178 279
rect 145 254 153 271
rect 170 254 178 271
rect 145 246 178 254
rect 212 271 245 279
rect 212 254 220 271
rect 237 254 245 271
rect 18 209 26 226
rect 43 225 51 226
rect 212 229 245 254
rect 212 225 220 229
rect 43 212 220 225
rect 237 212 245 229
rect 43 209 245 212
rect 18 208 245 209
rect 18 178 51 208
rect 18 161 26 178
rect 43 161 51 178
rect 18 153 51 161
rect 85 178 118 186
rect 85 161 93 178
rect 110 161 118 178
rect 85 153 118 161
rect 145 178 178 186
rect 145 161 153 178
rect 170 161 178 178
rect 145 153 178 161
rect 212 178 245 208
rect 212 161 220 178
rect 237 161 245 178
rect 212 153 245 161
rect 18 111 51 119
rect 18 94 26 111
rect 43 94 51 111
rect 18 86 51 94
rect 77 94 118 102
rect 77 77 93 94
rect 110 77 118 94
rect 77 70 118 77
rect 145 95 187 103
rect 145 78 153 95
rect 170 78 187 95
rect 145 70 187 78
rect 77 44 94 70
rect 170 61 187 70
rect 170 44 193 61
rect 11 9 44 17
rect 228 9 245 153
rect 0 -8 19 9
rect 36 -8 127 9
rect 144 -8 260 9
rect 11 -16 44 -8
<< viali >>
rect 36 504 53 521
rect 127 504 144 521
rect 140 358 157 375
rect 98 304 115 321
rect 26 94 43 111
rect 60 44 77 61
rect 193 44 210 61
rect 19 -8 36 9
rect 127 -8 144 9
<< metal1 >>
rect 0 526 260 527
rect 0 521 122 526
rect 0 504 36 521
rect 53 504 122 521
rect 0 500 122 504
rect 148 500 260 526
rect 0 498 260 500
rect 134 375 163 381
rect 134 358 140 375
rect 157 358 163 375
rect 134 352 163 358
rect 92 321 121 327
rect 92 304 98 321
rect 115 304 121 321
rect 92 298 121 304
rect 20 111 49 117
rect 20 101 26 111
rect 18 94 26 101
rect 43 101 49 111
rect 43 94 51 101
rect 18 86 51 94
rect 51 67 86 70
rect 51 38 54 67
rect 83 38 86 67
rect 51 35 86 38
rect 184 67 219 70
rect 184 38 187 67
rect 216 38 219 67
rect 184 35 219 38
rect 0 14 260 15
rect 0 9 122 14
rect 0 -8 19 9
rect 36 -8 122 9
rect 0 -12 122 -8
rect 148 -12 260 14
rect 0 -14 260 -12
<< via1 >>
rect 122 521 148 526
rect 122 504 127 521
rect 127 504 144 521
rect 144 504 148 521
rect 122 500 148 504
rect 54 61 83 67
rect 54 44 60 61
rect 60 44 77 61
rect 77 44 83 61
rect 54 38 83 44
rect 187 61 216 67
rect 187 44 193 61
rect 193 44 210 61
rect 210 44 216 61
rect 187 38 216 44
rect 122 9 148 14
rect 122 -8 127 9
rect 127 -8 144 9
rect 144 -8 148 9
rect 122 -12 148 -8
<< metal2 >>
rect 72 70 86 558
rect 113 529 156 534
rect 113 496 118 529
rect 151 496 156 529
rect 113 491 156 496
rect 51 67 86 70
rect 51 38 54 67
rect 83 38 86 67
rect 51 35 86 38
rect 72 -30 86 35
rect 184 70 198 560
rect 184 67 219 70
rect 184 38 187 67
rect 216 38 219 67
rect 184 35 219 38
rect 113 17 156 22
rect 113 -16 118 17
rect 151 -16 156 17
rect 113 -21 156 -16
rect 184 -30 198 35
<< via2 >>
rect 118 526 151 529
rect 118 500 122 526
rect 122 500 148 526
rect 148 500 151 526
rect 118 496 151 500
rect 118 14 151 17
rect 118 -12 122 14
rect 122 -12 148 14
rect 148 -12 151 14
rect 118 -16 151 -12
<< metal3 >>
rect 105 529 165 542
rect 105 496 118 529
rect 151 496 165 529
rect 105 482 165 496
rect 105 17 165 30
rect 105 -16 118 17
rect 151 -16 165 17
rect 105 -30 165 -16
<< labels >>
flabel metal1 s 28 96 41 107 0 FreeSans 200 0 0 0 wl
port 3 nsew
flabel metal1 s 38 509 51 520 0 FreeSans 200 0 0 0 vdd
port 4 nsew
flabel metal1 s 143 361 154 372 0 FreeSans 200 0 0 0 Q_bar
flabel metal1 s 102 308 113 319 0 FreeSans 200 0 0 0 Q
flabel metal1 s 22 -4 35 7 0 FreeSans 200 0 0 0 gnd
port 5 nsew
flabel metal2 s 74 20 83 31 0 FreeSans 200 0 0 0 bl
port 0 nsew
flabel metal2 s 187 21 196 32 0 FreeSans 200 0 0 0 br
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 260 513
<< end >>
