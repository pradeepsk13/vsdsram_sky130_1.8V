magic
tech sky130A
timestamp 1605371449
<< nwell >>
rect 511 334 837 529
<< nmos >>
rect 600 76 615 202
rect 740 75 755 201
rect 620 -82 662 -67
rect 758 -82 800 -67
<< pmos >>
rect 600 364 615 419
rect 740 364 755 419
<< ndiff >>
rect 555 161 600 202
rect 555 144 568 161
rect 585 144 600 161
rect 555 108 600 144
rect 555 91 568 108
rect 585 91 600 108
rect 555 76 600 91
rect 615 161 660 202
rect 615 144 628 161
rect 645 144 660 161
rect 615 108 660 144
rect 615 91 628 108
rect 645 91 660 108
rect 615 76 660 91
rect 700 160 740 201
rect 700 143 708 160
rect 725 143 740 160
rect 700 107 740 143
rect 700 90 708 107
rect 725 90 740 107
rect 700 75 740 90
rect 755 160 800 201
rect 755 143 768 160
rect 785 143 800 160
rect 755 107 800 143
rect 755 90 768 107
rect 785 90 800 107
rect 755 75 800 90
rect 620 -37 662 -27
rect 620 -54 633 -37
rect 650 -54 662 -37
rect 620 -67 662 -54
rect 758 -37 800 -27
rect 758 -54 771 -37
rect 788 -54 800 -37
rect 758 -67 800 -54
rect 620 -95 662 -82
rect 620 -112 633 -95
rect 650 -112 662 -95
rect 620 -127 662 -112
rect 758 -95 800 -82
rect 758 -112 771 -95
rect 788 -112 800 -95
rect 758 -127 800 -112
<< pdiff >>
rect 558 401 600 419
rect 558 384 568 401
rect 585 384 600 401
rect 558 364 600 384
rect 615 401 660 419
rect 615 384 628 401
rect 645 384 660 401
rect 615 364 660 384
rect 698 401 740 419
rect 698 384 708 401
rect 725 384 740 401
rect 698 364 740 384
rect 755 401 800 419
rect 755 384 768 401
rect 785 384 800 401
rect 755 364 800 384
<< ndiffc >>
rect 568 144 585 161
rect 568 91 585 108
rect 628 144 645 161
rect 628 91 645 108
rect 708 143 725 160
rect 708 90 725 107
rect 768 143 785 160
rect 768 90 785 107
rect 633 -54 650 -37
rect 771 -54 788 -37
rect 633 -112 650 -95
rect 771 -112 788 -95
<< pdiffc >>
rect 568 384 585 401
rect 628 384 645 401
rect 708 384 725 401
rect 768 384 785 401
<< psubdiff >>
rect 563 -190 604 -178
rect 563 -207 575 -190
rect 592 -207 604 -190
rect 563 -219 604 -207
rect 691 -190 732 -178
rect 691 -207 703 -190
rect 720 -207 732 -190
rect 691 -219 732 -207
rect 804 -190 845 -178
rect 804 -207 816 -190
rect 833 -207 845 -190
rect 804 -219 845 -207
<< nsubdiff >>
rect 562 495 595 496
rect 562 484 685 495
rect 562 467 574 484
rect 591 467 685 484
rect 562 455 685 467
rect 771 483 812 495
rect 771 466 783 483
rect 800 466 812 483
rect 771 454 812 466
<< psubdiffcont >>
rect 575 -207 592 -190
rect 703 -207 720 -190
rect 816 -207 833 -190
<< nsubdiffcont >>
rect 574 467 591 484
rect 783 466 800 483
<< poly >>
rect 600 419 615 434
rect 740 419 755 434
rect 600 270 615 364
rect 740 333 755 364
rect 722 325 755 333
rect 722 308 730 325
rect 747 308 755 325
rect 722 300 755 308
rect 582 262 615 270
rect 582 245 590 262
rect 607 245 615 262
rect 582 237 615 245
rect 600 202 615 237
rect 740 201 755 300
rect 600 60 615 76
rect 740 60 755 75
rect 548 -65 583 -56
rect 548 -82 557 -65
rect 574 -67 583 -65
rect 574 -82 620 -67
rect 662 -82 758 -67
rect 800 -82 820 -67
rect 548 -91 583 -82
<< polycont >>
rect 730 308 747 325
rect 590 245 607 262
rect 557 -82 574 -65
<< locali >>
rect 485 495 595 496
rect 485 484 882 495
rect 485 467 544 484
rect 561 467 574 484
rect 591 483 882 484
rect 591 467 730 483
rect 485 466 730 467
rect 747 466 783 483
rect 800 466 817 483
rect 834 466 882 483
rect 485 455 882 466
rect 565 409 585 455
rect 705 409 725 455
rect 560 401 593 409
rect 560 384 568 401
rect 585 384 593 401
rect 560 376 593 384
rect 620 401 653 409
rect 620 384 628 401
rect 645 384 653 401
rect 620 376 653 384
rect 700 401 733 409
rect 700 384 708 401
rect 725 384 733 401
rect 700 376 733 384
rect 760 401 793 409
rect 760 384 768 401
rect 785 384 793 401
rect 760 376 793 384
rect 635 325 653 376
rect 722 325 755 333
rect 635 308 730 325
rect 747 308 755 325
rect 635 305 755 308
rect 582 262 615 270
rect 582 245 590 262
rect 607 245 615 262
rect 582 237 615 245
rect 635 202 653 305
rect 722 300 755 305
rect 775 266 793 376
rect 769 260 798 266
rect 769 243 775 260
rect 792 243 798 260
rect 769 237 798 243
rect 560 161 593 202
rect 560 144 568 161
rect 585 144 593 161
rect 560 108 593 144
rect 560 91 568 108
rect 585 91 593 108
rect 560 83 593 91
rect 620 161 653 202
rect 775 201 793 237
rect 620 144 628 161
rect 645 144 653 161
rect 620 108 653 144
rect 620 91 628 108
rect 645 91 653 108
rect 620 83 653 91
rect 700 160 733 201
rect 700 143 708 160
rect 725 143 733 160
rect 700 107 733 143
rect 700 90 708 107
rect 725 90 733 107
rect 570 23 590 83
rect 561 17 590 23
rect 561 0 567 17
rect 584 0 590 17
rect 561 -6 590 0
rect 625 -29 645 83
rect 700 82 733 90
rect 760 160 793 201
rect 760 143 768 160
rect 785 143 793 160
rect 760 107 793 143
rect 760 90 768 107
rect 785 90 793 107
rect 760 82 793 90
rect 710 23 730 82
rect 701 17 730 23
rect 701 0 707 17
rect 724 0 730 17
rect 701 -6 730 0
rect 625 -37 658 -29
rect 625 -54 633 -37
rect 650 -54 658 -37
rect 548 -65 583 -56
rect 625 -62 658 -54
rect 548 -82 557 -65
rect 574 -82 583 -65
rect 548 -91 583 -82
rect 625 -95 658 -87
rect 625 -112 633 -95
rect 650 -112 658 -95
rect 625 -120 658 -112
rect 548 -131 577 -125
rect 548 -148 554 -131
rect 571 -134 577 -131
rect 625 -134 645 -120
rect 571 -148 645 -134
rect 548 -154 645 -148
rect 705 -182 725 -6
rect 772 -29 792 82
rect 763 -37 796 -29
rect 763 -54 771 -37
rect 788 -54 796 -37
rect 763 -62 796 -54
rect 763 -95 796 -87
rect 763 -112 771 -95
rect 788 -112 796 -95
rect 763 -120 796 -112
rect 775 -139 795 -120
rect 841 -136 870 -130
rect 841 -139 847 -136
rect 775 -153 847 -139
rect 864 -153 870 -136
rect 775 -159 870 -153
rect 567 -190 841 -182
rect 567 -207 575 -190
rect 592 -207 638 -190
rect 655 -207 703 -190
rect 720 -207 759 -190
rect 776 -207 816 -190
rect 833 -207 841 -190
rect 567 -215 841 -207
<< viali >>
rect 544 467 561 484
rect 730 466 747 483
rect 817 466 834 483
rect 590 245 607 262
rect 775 243 792 260
rect 567 0 584 17
rect 707 0 724 17
rect 554 -148 571 -131
rect 847 -153 864 -136
rect 638 -207 655 -190
rect 759 -207 776 -190
<< metal1 >>
rect 485 495 595 496
rect 485 484 882 495
rect 485 467 544 484
rect 561 483 882 484
rect 561 467 730 483
rect 485 466 730 467
rect 747 466 817 483
rect 834 466 882 483
rect 485 455 882 466
rect 582 262 615 270
rect 582 245 590 262
rect 607 260 615 262
rect 769 260 798 266
rect 607 245 775 260
rect 582 243 775 245
rect 792 243 798 260
rect 582 240 798 243
rect 582 237 615 240
rect 769 237 798 240
rect 561 20 590 23
rect 701 20 730 23
rect 561 17 730 20
rect 561 0 567 17
rect 584 0 707 17
rect 724 0 730 17
rect 561 -6 590 0
rect 701 -6 730 0
rect 548 -131 577 -125
rect 548 -148 554 -131
rect 571 -148 577 -131
rect 548 -154 577 -148
rect 841 -136 870 -130
rect 841 -153 847 -136
rect 864 -153 870 -136
rect 841 -159 870 -153
rect 548 -190 850 -175
rect 548 -207 638 -190
rect 655 -207 759 -190
rect 776 -207 850 -190
rect 548 -219 850 -207
<< labels >>
flabel metal1 s 494 463 537 488 0 FreeSans 240 0 0 0 vdd
port 1 nsew
flabel locali s 733 310 742 321 0 FreeSans 200 0 0 0 q
port 6 nsew
flabel locali s 591 247 602 257 0 FreeSans 200 0 0 0 qb
port 7 nsew
flabel metal1 s 661 -209 704 -184 0 FreeSans 240 0 0 0 gnd
port 2 nsew
flabel locali s 558 -81 566 -69 0 FreeSans 240 0 0 0 wl
port 3 nsew
flabel locali s 557 -146 565 -134 0 FreeSans 240 0 0 0 bl
port 4 nsew
flabel locali s 849 -149 857 -137 0 FreeSans 240 0 0 0 blb
port 5 nsew
<< end >>
