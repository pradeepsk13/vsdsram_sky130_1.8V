magic
tech sky130A
timestamp 1616270591
<< nwell >>
rect 0 273 1271 453
<< nmos >>
rect 64 57 79 99
rect 207 57 222 99
rect 328 57 343 99
rect 499 57 514 99
rect 594 57 609 99
rect 787 57 802 99
rect 908 57 923 99
rect 1103 57 1118 99
rect 1198 57 1213 99
<< pmos >>
rect 64 291 79 346
rect 207 291 222 346
rect 328 291 343 346
rect 499 291 514 346
rect 594 291 609 346
rect 787 291 802 346
rect 908 291 923 346
rect 1103 291 1118 346
rect 1198 291 1213 346
<< ndiff >>
rect 18 88 64 99
rect 18 71 28 88
rect 45 71 64 88
rect 18 57 64 71
rect 79 88 125 99
rect 79 71 97 88
rect 114 71 125 88
rect 79 57 125 71
rect 161 88 207 99
rect 161 71 171 88
rect 188 71 207 88
rect 161 57 207 71
rect 222 88 328 99
rect 222 71 281 88
rect 298 71 328 88
rect 222 57 328 71
rect 343 88 411 99
rect 343 71 376 88
rect 393 71 411 88
rect 343 57 411 71
rect 446 87 499 99
rect 446 70 459 87
rect 476 70 499 87
rect 446 57 499 70
rect 514 88 594 99
rect 514 71 547 88
rect 564 71 594 88
rect 514 57 594 71
rect 609 88 671 99
rect 609 71 622 88
rect 639 71 671 88
rect 609 57 671 71
rect 722 88 787 99
rect 722 71 751 88
rect 768 71 787 88
rect 722 57 787 71
rect 802 88 908 99
rect 802 71 861 88
rect 878 71 908 88
rect 802 57 908 71
rect 923 88 1002 99
rect 923 71 956 88
rect 973 71 1002 88
rect 923 57 1002 71
rect 1047 88 1103 99
rect 1047 71 1063 88
rect 1080 71 1103 88
rect 1047 57 1103 71
rect 1118 88 1198 99
rect 1118 71 1151 88
rect 1168 71 1198 88
rect 1118 57 1198 71
rect 1213 88 1253 99
rect 1213 71 1226 88
rect 1243 71 1253 88
rect 1213 57 1253 71
<< pdiff >>
rect 18 328 64 346
rect 18 311 28 328
rect 45 311 64 328
rect 18 291 64 311
rect 79 328 125 346
rect 79 311 97 328
rect 114 311 125 328
rect 79 291 125 311
rect 161 328 207 346
rect 161 311 171 328
rect 188 311 207 328
rect 161 291 207 311
rect 222 328 328 346
rect 222 311 281 328
rect 298 311 328 328
rect 222 291 328 311
rect 343 328 411 346
rect 343 311 376 328
rect 393 311 411 328
rect 343 291 411 311
rect 446 328 499 346
rect 446 311 464 328
rect 481 311 499 328
rect 446 291 499 311
rect 514 328 594 346
rect 514 311 547 328
rect 564 311 594 328
rect 514 291 594 311
rect 609 328 672 346
rect 609 311 622 328
rect 639 311 672 328
rect 609 291 672 311
rect 723 328 787 346
rect 723 311 751 328
rect 768 311 787 328
rect 723 291 787 311
rect 802 328 908 346
rect 802 311 861 328
rect 878 311 908 328
rect 802 291 908 311
rect 923 328 1002 346
rect 923 311 956 328
rect 973 311 1002 328
rect 923 291 1002 311
rect 1047 328 1103 346
rect 1047 311 1060 328
rect 1077 311 1103 328
rect 1047 291 1103 311
rect 1118 328 1198 346
rect 1118 311 1151 328
rect 1168 311 1198 328
rect 1118 291 1198 311
rect 1213 328 1253 346
rect 1213 311 1226 328
rect 1243 311 1253 328
rect 1213 291 1253 311
<< ndiffc >>
rect 28 71 45 88
rect 97 71 114 88
rect 171 71 188 88
rect 281 71 298 88
rect 376 71 393 88
rect 459 70 476 87
rect 547 71 564 88
rect 622 71 639 88
rect 751 71 768 88
rect 861 71 878 88
rect 956 71 973 88
rect 1063 71 1080 88
rect 1151 71 1168 88
rect 1226 71 1243 88
<< pdiffc >>
rect 28 311 45 328
rect 97 311 114 328
rect 171 311 188 328
rect 281 311 298 328
rect 376 311 393 328
rect 464 311 481 328
rect 547 311 564 328
rect 622 311 639 328
rect 751 311 768 328
rect 861 311 878 328
rect 956 311 973 328
rect 1060 311 1077 328
rect 1151 311 1168 328
rect 1226 311 1243 328
<< psubdiff >>
rect 3 8 44 20
rect 3 -9 15 8
rect 32 -9 44 8
rect 3 -21 44 -9
rect 146 8 187 20
rect 146 -9 158 8
rect 175 -9 187 8
rect 146 -21 187 -9
rect 250 8 291 20
rect 250 -9 262 8
rect 279 -9 291 8
rect 250 -21 291 -9
rect 361 8 402 20
rect 361 -9 373 8
rect 390 -9 402 8
rect 361 -21 402 -9
rect 546 8 587 20
rect 546 -9 558 8
rect 575 -9 587 8
rect 546 -21 587 -9
rect 726 8 767 20
rect 726 -9 738 8
rect 755 -9 767 8
rect 726 -21 767 -9
rect 830 8 871 20
rect 830 -9 842 8
rect 859 -9 871 8
rect 830 -21 871 -9
rect 941 8 982 20
rect 941 -9 953 8
rect 970 -9 982 8
rect 941 -21 982 -9
rect 1150 8 1191 20
rect 1150 -9 1162 8
rect 1179 -9 1191 8
rect 1150 -21 1191 -9
<< nsubdiff >>
rect 18 417 71 435
rect 18 400 36 417
rect 53 400 71 417
rect 18 382 71 400
rect 161 417 214 435
rect 161 400 179 417
rect 196 400 214 417
rect 161 382 214 400
rect 313 417 366 435
rect 313 400 331 417
rect 348 400 366 417
rect 313 382 366 400
rect 547 417 600 435
rect 547 400 565 417
rect 582 400 600 417
rect 547 382 600 400
rect 741 417 794 435
rect 741 400 759 417
rect 776 400 794 417
rect 741 382 794 400
rect 893 417 946 435
rect 893 400 911 417
rect 928 400 946 417
rect 893 382 946 400
rect 1151 417 1204 435
rect 1151 400 1169 417
rect 1186 400 1204 417
rect 1151 382 1204 400
<< psubdiffcont >>
rect 15 -9 32 8
rect 158 -9 175 8
rect 262 -9 279 8
rect 373 -9 390 8
rect 558 -9 575 8
rect 738 -9 755 8
rect 842 -9 859 8
rect 953 -9 970 8
rect 1162 -9 1179 8
<< nsubdiffcont >>
rect 36 400 53 417
rect 179 400 196 417
rect 331 400 348 417
rect 565 400 582 417
rect 759 400 776 417
rect 911 400 928 417
rect 1169 400 1186 417
<< poly >>
rect 64 346 79 361
rect 207 346 222 361
rect 328 346 343 361
rect 499 346 514 361
rect 594 346 609 361
rect 787 346 802 361
rect 908 346 923 361
rect 1103 346 1118 361
rect 1198 346 1213 361
rect 8 218 41 226
rect 8 201 16 218
rect 33 217 41 218
rect 64 219 79 291
rect 207 219 222 291
rect 328 269 343 291
rect 499 271 514 291
rect 319 261 352 269
rect 319 244 327 261
rect 344 244 352 261
rect 319 236 352 244
rect 499 263 532 271
rect 499 246 507 263
rect 524 246 532 263
rect 499 238 532 246
rect 64 217 222 219
rect 33 215 222 217
rect 33 207 352 215
rect 33 202 327 207
rect 33 201 41 202
rect 8 193 41 201
rect 64 199 327 202
rect 64 99 79 199
rect 319 190 327 199
rect 344 190 352 207
rect 319 182 352 190
rect 207 162 240 170
rect 207 145 215 162
rect 232 145 240 162
rect 207 137 240 145
rect 207 99 222 137
rect 328 99 343 182
rect 499 99 514 238
rect 594 154 609 291
rect 727 262 760 269
rect 787 262 802 291
rect 908 269 923 291
rect 727 261 802 262
rect 727 244 735 261
rect 752 247 802 261
rect 752 244 760 247
rect 727 236 760 244
rect 787 215 802 247
rect 899 261 932 269
rect 899 244 907 261
rect 924 244 932 261
rect 899 236 932 244
rect 1103 234 1118 291
rect 1103 226 1136 234
rect 787 207 932 215
rect 787 199 907 207
rect 899 190 907 199
rect 924 190 932 207
rect 899 182 932 190
rect 1103 209 1111 226
rect 1128 209 1136 226
rect 1103 201 1136 209
rect 576 146 609 154
rect 576 129 584 146
rect 601 129 609 146
rect 576 121 609 129
rect 594 99 609 121
rect 787 162 820 170
rect 787 145 795 162
rect 812 145 820 162
rect 787 137 820 145
rect 787 99 802 137
rect 908 99 923 182
rect 1103 99 1118 201
rect 1198 150 1213 291
rect 1180 142 1213 150
rect 1180 125 1188 142
rect 1205 125 1213 142
rect 1180 117 1213 125
rect 1198 99 1213 117
rect 64 42 79 57
rect 207 42 222 57
rect 328 42 343 57
rect 499 42 514 57
rect 594 42 609 57
rect 787 42 802 57
rect 908 42 923 57
rect 1103 42 1118 57
rect 1198 42 1213 57
<< polycont >>
rect 16 201 33 218
rect 327 244 344 261
rect 507 246 524 263
rect 327 190 344 207
rect 215 145 232 162
rect 735 244 752 261
rect 907 244 924 261
rect 907 190 924 207
rect 1111 209 1128 226
rect 584 129 601 146
rect 795 145 812 162
rect 1188 125 1205 142
<< locali >>
rect 6 417 1271 425
rect 6 400 36 417
rect 53 400 179 417
rect 196 400 258 417
rect 275 400 331 417
rect 348 400 486 417
rect 503 400 565 417
rect 582 400 644 417
rect 661 400 759 417
rect 776 400 838 417
rect 855 400 911 417
rect 928 400 1090 417
rect 1107 400 1169 417
rect 1186 400 1248 417
rect 1265 400 1271 417
rect 6 392 1271 400
rect 26 336 46 392
rect 542 336 562 392
rect 1146 336 1166 392
rect 20 328 53 336
rect 20 311 28 328
rect 45 311 53 328
rect 20 303 53 311
rect 89 328 122 336
rect 89 311 97 328
rect 114 311 122 328
rect 89 303 122 311
rect 163 328 196 336
rect 163 311 171 328
rect 188 311 196 328
rect 163 303 196 311
rect 273 328 306 336
rect 273 311 281 328
rect 298 311 306 328
rect 273 303 306 311
rect 368 332 401 336
rect 456 332 489 336
rect 368 328 489 332
rect 368 311 376 328
rect 393 311 464 328
rect 481 311 489 328
rect 368 307 489 311
rect 368 303 401 307
rect 456 303 489 307
rect 539 328 572 336
rect 539 311 547 328
rect 564 311 572 328
rect 539 303 572 311
rect 614 328 776 336
rect 614 311 622 328
rect 639 311 751 328
rect 768 311 776 328
rect 614 303 776 311
rect 853 328 886 336
rect 853 311 861 328
rect 878 311 886 328
rect 853 303 886 311
rect 948 328 981 336
rect 948 311 956 328
rect 973 327 981 328
rect 1052 328 1085 336
rect 1052 327 1060 328
rect 973 311 1060 327
rect 1077 311 1085 328
rect 948 307 1085 311
rect 948 303 981 307
rect 1052 303 1085 307
rect 1143 328 1176 336
rect 1143 311 1151 328
rect 1168 311 1176 328
rect 1143 303 1176 311
rect 1218 328 1251 336
rect 1218 311 1226 328
rect 1243 311 1251 328
rect 1218 303 1251 311
rect 8 218 41 226
rect 8 201 16 218
rect 33 201 41 218
rect 8 175 41 201
rect 8 158 16 175
rect 33 158 41 175
rect 96 168 116 303
rect 166 263 186 303
rect 158 257 186 263
rect 158 240 163 257
rect 180 240 186 257
rect 158 235 186 240
rect 8 151 41 158
rect 95 162 124 168
rect 95 145 101 162
rect 118 145 124 162
rect 95 139 124 145
rect 96 96 116 139
rect 166 96 186 235
rect 207 162 240 170
rect 207 145 215 162
rect 232 145 240 162
rect 207 137 240 145
rect 278 157 298 303
rect 319 261 352 269
rect 319 244 327 261
rect 344 244 352 261
rect 319 236 352 244
rect 319 207 352 215
rect 319 190 327 207
rect 344 190 352 207
rect 319 182 352 190
rect 278 149 310 157
rect 278 132 286 149
rect 303 132 310 149
rect 278 126 310 132
rect 278 96 298 126
rect 373 96 393 303
rect 499 264 532 271
rect 627 264 647 303
rect 499 263 647 264
rect 499 246 507 263
rect 524 246 647 263
rect 499 244 647 246
rect 499 238 532 244
rect 576 146 609 154
rect 576 129 584 146
rect 601 129 609 146
rect 576 121 609 129
rect 627 96 647 244
rect 727 261 760 269
rect 727 244 735 261
rect 752 244 760 261
rect 727 236 760 244
rect 787 162 820 170
rect 787 145 795 162
rect 812 145 820 162
rect 787 137 820 145
rect 858 158 878 303
rect 899 261 932 269
rect 899 244 907 261
rect 924 244 932 261
rect 899 236 932 244
rect 899 207 932 215
rect 899 190 907 207
rect 924 190 932 207
rect 899 182 932 190
rect 858 150 890 158
rect 858 133 866 150
rect 883 133 890 150
rect 858 127 890 133
rect 858 96 878 127
rect 953 96 973 303
rect 1045 227 1136 234
rect 1231 227 1251 303
rect 1045 226 1251 227
rect 1045 209 1052 226
rect 1069 209 1111 226
rect 1128 209 1251 226
rect 1045 207 1251 209
rect 1045 202 1136 207
rect 1103 201 1136 202
rect 1180 142 1213 150
rect 1180 125 1188 142
rect 1205 125 1213 142
rect 1180 117 1213 125
rect 1231 96 1251 207
rect 20 88 53 96
rect 20 71 28 88
rect 45 71 53 88
rect 20 63 53 71
rect 89 88 122 96
rect 89 71 97 88
rect 114 71 122 88
rect 89 63 122 71
rect 163 88 196 96
rect 163 71 171 88
rect 188 71 196 88
rect 163 63 196 71
rect 273 88 306 96
rect 273 71 281 88
rect 298 71 306 88
rect 273 63 306 71
rect 368 88 401 96
rect 368 71 376 88
rect 393 87 401 88
rect 451 87 484 95
rect 393 71 459 87
rect 368 70 459 71
rect 476 70 484 87
rect 368 67 484 70
rect 368 63 401 67
rect 26 16 46 63
rect 451 62 484 67
rect 539 88 572 96
rect 539 71 547 88
rect 564 71 572 88
rect 539 63 572 71
rect 552 16 572 63
rect 614 88 776 96
rect 614 71 622 88
rect 639 71 751 88
rect 768 71 776 88
rect 614 62 776 71
rect 853 88 886 96
rect 853 71 861 88
rect 878 71 886 88
rect 853 63 886 71
rect 948 88 981 96
rect 948 71 956 88
rect 973 87 981 88
rect 1055 88 1088 96
rect 1055 87 1063 88
rect 973 71 1063 87
rect 1080 71 1088 88
rect 948 67 1088 71
rect 948 63 981 67
rect 1055 63 1088 67
rect 1143 88 1176 96
rect 1143 71 1151 88
rect 1168 71 1176 88
rect 1143 63 1176 71
rect 1218 88 1251 96
rect 1218 71 1226 88
rect 1243 71 1251 88
rect 1218 63 1251 71
rect 1156 16 1176 63
rect 0 8 1253 16
rect 0 -9 15 8
rect 32 -9 75 8
rect 92 -9 158 8
rect 175 -9 218 8
rect 235 -9 262 8
rect 279 -9 322 8
rect 339 -9 373 8
rect 390 -9 509 8
rect 526 -9 558 8
rect 575 -9 618 8
rect 635 -9 738 8
rect 755 -9 798 8
rect 815 -9 842 8
rect 859 -9 902 8
rect 919 -9 953 8
rect 970 -9 1113 8
rect 1130 -9 1162 8
rect 1179 -9 1222 8
rect 1239 -9 1253 8
rect 0 -17 1253 -9
<< viali >>
rect 258 400 275 417
rect 486 400 503 417
rect 644 400 661 417
rect 838 400 855 417
rect 1090 400 1107 417
rect 1248 400 1265 417
rect 16 158 33 175
rect 163 240 180 257
rect 101 145 118 162
rect 215 145 232 162
rect 327 244 344 261
rect 327 190 344 207
rect 286 132 303 149
rect 584 129 601 146
rect 735 244 752 261
rect 795 145 812 162
rect 907 244 924 261
rect 866 133 883 150
rect 1052 209 1069 226
rect 1188 125 1205 142
rect 75 -9 92 8
rect 218 -9 235 8
rect 322 -9 339 8
rect 509 -9 526 8
rect 618 -9 635 8
rect 798 -9 815 8
rect 902 -9 919 8
rect 1113 -9 1130 8
rect 1222 -9 1239 8
<< metal1 >>
rect 6 417 1271 425
rect 6 400 258 417
rect 275 400 486 417
rect 503 400 644 417
rect 661 400 838 417
rect 855 400 1090 417
rect 1107 400 1248 417
rect 1265 400 1271 417
rect 6 392 1271 400
rect 123 262 186 265
rect 123 236 127 262
rect 153 257 186 262
rect 319 261 352 269
rect 319 257 327 261
rect 153 240 163 257
rect 180 240 186 257
rect 153 236 186 240
rect 123 233 186 236
rect 211 244 327 257
rect 344 257 352 261
rect 727 261 760 269
rect 727 257 735 261
rect 344 244 735 257
rect 752 244 760 261
rect 899 261 932 269
rect 899 257 907 261
rect 211 237 760 244
rect 8 180 76 183
rect 8 175 47 180
rect 8 158 16 175
rect 33 158 47 175
rect 8 154 47 158
rect 73 154 76 180
rect 211 170 231 237
rect 319 236 352 237
rect 727 236 760 237
rect 791 244 907 257
rect 924 244 932 261
rect 791 237 932 244
rect 319 212 352 215
rect 791 212 811 237
rect 899 236 932 237
rect 319 207 811 212
rect 319 190 327 207
rect 344 190 811 207
rect 1013 231 1076 234
rect 1013 205 1016 231
rect 1042 226 1076 231
rect 1042 209 1052 226
rect 1069 209 1076 226
rect 1042 205 1076 209
rect 1013 202 1076 205
rect 319 187 811 190
rect 319 182 352 187
rect 791 170 811 187
rect 8 151 76 154
rect 95 162 124 168
rect 207 162 240 170
rect 95 145 101 162
rect 118 145 215 162
rect 232 145 240 162
rect 787 162 820 170
rect 95 142 240 145
rect 95 139 124 142
rect 207 137 240 142
rect 280 149 310 157
rect 280 132 286 149
rect 303 147 310 149
rect 576 147 609 154
rect 303 146 609 147
rect 303 132 584 146
rect 280 129 584 132
rect 601 129 609 146
rect 787 145 795 162
rect 812 145 820 162
rect 787 137 820 145
rect 860 150 890 158
rect 280 126 609 129
rect 860 133 866 150
rect 883 147 890 150
rect 1179 147 1213 150
rect 883 142 1213 147
rect 883 133 1188 142
rect 860 127 1188 133
rect 576 121 609 126
rect 1179 125 1188 127
rect 1205 125 1213 142
rect 1179 117 1213 125
rect 0 8 1253 16
rect 0 -9 75 8
rect 92 -9 218 8
rect 235 -9 322 8
rect 339 -9 509 8
rect 526 -9 618 8
rect 635 -9 798 8
rect 815 -9 902 8
rect 919 -9 1113 8
rect 1130 -9 1222 8
rect 1239 -9 1253 8
rect 0 -17 1253 -9
<< via1 >>
rect 127 236 153 262
rect 47 154 73 180
rect 1016 205 1042 231
<< metal2 >>
rect 123 262 157 265
rect 123 236 127 262
rect 153 236 157 262
rect 123 233 157 236
rect 1013 231 1045 234
rect 1013 205 1016 231
rect 1042 205 1045 231
rect 1013 202 1045 205
rect 45 180 76 183
rect 45 154 47 180
rect 73 154 76 180
rect 45 151 76 154
<< labels >>
flabel metal2 s 127 236 153 262 0 FreeSans 400 0 0 0 D
port 0 nsew
flabel locali s 289 136 297 143 0 FreeSans 200 0 0 0 net1
flabel locali s 379 162 387 170 0 FreeSans 200 0 0 0 net2
flabel metal1 s 539 -17 674 16 0 FreeSans 400 0 0 0 gnd
port 4 nsew
flabel locali s 635 130 643 138 0 FreeSans 200 0 0 0 net3
flabel locali s 871 136 879 143 0 FreeSans 200 0 0 0 net4
flabel locali s 958 312 968 324 0 FreeSans 200 0 0 0 net5
flabel locali s 217 146 228 159 0 FreeSans 240 0 0 0 clkb
flabel metal2 s 1016 205 1042 231 0 FreeSans 400 0 0 0 Q
port 1 nsew
flabel metal2 s 47 154 73 180 0 FreeSans 200 0 0 0 clk
port 2 nsew
flabel metal1 s 592 398 631 418 0 FreeSans 400 0 0 0 vdd
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1271 409
<< end >>
