* NGSPICE file created from sram_ip.ext - technology: sky130A

.subckt sram_ip din wb gnd vdd blb bl qb q wl rd_en dout
X0 net7 net6 vdd vdd sky130_fd_pr__pfet_01v8 w=1e+06u l=150000u
X1 net2 wb net3 vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X2 q qb gnd gnd sky130_fd_pr__nfet_01v8 w=1.26e+06u l=150000u
X3 qb wl blb gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 bl gnd vdd vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X5 net3 net1 vdd vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X6 q wl bl gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 bl net5 gnd gnd sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 net5 wb net9 vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X9 q qb vdd vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X10 dout net7 vdd vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X11 blb net2 gnd gnd sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 net1 din vdd vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X13 qb q vdd vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X14 net7 bl net8 gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 net5 net4 gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 net8 rd_en gnd gnd sky130_fd_pr__nfet_01v8 w=1e+06u l=150000u
X17 vdd net6 net6 vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X18 net8 blb net6 gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 blb gnd vdd vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X20 net1 din gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 net9 net4 vdd vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
X22 net2 net1 gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 net2 wb gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 net4 net1 gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 qb q gnd gnd sky130_fd_pr__nfet_01v8 w=1.26e+06u l=150000u
X26 dout net7 gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 net5 wb gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 net4 net1 vdd vdd sky130_fd_pr__pfet_01v8 w=550000u l=150000u
C0 net7 net6 0.09fF
C1 net3 blb 0.02fF
C2 net2 net1 0.09fF
C3 net3 vdd 0.29fF
C4 blb bl 0.58fF
C5 net4 net1 0.04fF
C6 q blb 0.22fF
C7 net2 wb 0.04fF
C8 qb bl 0.04fF
C9 net8 bl 0.06fF
C10 net9 vdd 0.27fF
C11 bl vdd 0.26fF
C12 wl bl 0.07fF
C13 net6 bl 0.01fF
C14 net5 vdd 0.06fF
C15 qb q 0.43fF
C16 q vdd 0.32fF
C17 wl q 0.01fF
C18 net7 bl 0.03fF
C19 net4 wb 0.05fF
C20 net6 q 0.09fF
C21 rd_en dout 0.01fF
C22 net1 vdd 0.41fF
C23 din vdd 0.07fF
C24 wb vdd 0.04fF
C25 net9 net5 0.21fF
C26 net5 bl 0.14fF
C27 q bl 0.30fF
C28 net3 net1 0.04fF
C29 dout vdd 0.15fF
C30 net2 blb 0.15fF
C31 net7 dout 0.09fF
C32 net2 vdd 0.21fF
C33 rd_en qb 0.01fF
C34 net8 rd_en 0.01fF
C35 rd_en vdd 0.03fF
C36 net9 wb 0.05fF
C37 wb bl 0.01fF
C38 net6 rd_en 0.02fF
C39 net4 vdd 0.32fF
C40 net5 wb 0.15fF
C41 net7 rd_en 0.01fF
C42 net3 net2 0.22fF
C43 net1 din 0.06fF
C44 qb blb 0.21fF
C45 net8 blb 0.02fF
C46 blb vdd 0.28fF
C47 net1 wb 0.05fF
C48 wl blb 0.12fF
C49 net6 blb 0.05fF
C50 net2 bl 0.01fF
C51 net8 qb 0.01fF
C52 qb vdd 0.37fF
C53 net8 vdd 0.00fF
C54 wl qb 0.01fF
C55 net6 qb 0.20fF
C56 net6 net8 0.19fF
C57 net6 vdd 0.34fF
C58 net4 net9 0.04fF
C59 net7 net8 0.25fF
C60 net7 vdd 0.26fF
C61 net4 net5 0.08fF
.ends

