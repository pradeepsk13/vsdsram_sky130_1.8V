magic
tech sky130A
timestamp 1616958208
<< nwell >>
rect 0 283 308 468
<< nmos >>
rect 250 199 265 241
rect 90 176 216 191
rect 90 126 216 141
rect 250 76 265 118
<< pmos >>
rect 101 302 116 357
rect 214 302 229 357
<< ndiff >>
rect 90 233 250 241
rect 90 216 98 233
rect 115 216 144 233
rect 161 216 179 233
rect 196 216 250 233
rect 90 199 250 216
rect 265 233 299 241
rect 265 216 274 233
rect 291 216 299 233
rect 265 199 299 216
rect 90 191 216 199
rect 90 167 216 176
rect 90 150 98 167
rect 115 150 141 167
rect 158 150 179 167
rect 196 150 216 167
rect 90 141 216 150
rect 90 118 216 126
rect 90 101 250 118
rect 90 84 98 101
rect 115 84 224 101
rect 241 84 250 101
rect 90 76 250 84
rect 265 101 299 118
rect 265 84 275 101
rect 292 84 299 101
rect 265 76 299 84
<< pdiff >>
rect 66 349 101 357
rect 66 332 74 349
rect 91 332 101 349
rect 66 302 101 332
rect 116 327 151 357
rect 116 310 126 327
rect 143 310 151 327
rect 116 302 151 310
rect 179 349 214 357
rect 179 332 187 349
rect 204 332 214 349
rect 179 302 214 332
rect 229 327 264 357
rect 229 310 239 327
rect 256 310 264 327
rect 229 302 264 310
<< ndiffc >>
rect 98 216 115 233
rect 144 216 161 233
rect 179 216 196 233
rect 274 216 291 233
rect 98 150 115 167
rect 141 150 158 167
rect 179 150 196 167
rect 98 84 115 101
rect 224 84 241 101
rect 275 84 292 101
<< pdiffc >>
rect 74 332 91 349
rect 126 310 143 327
rect 187 332 204 349
rect 239 310 256 327
<< psubdiff >>
rect 42 9 83 21
rect 42 -8 54 9
rect 71 -8 83 9
rect 42 -20 83 -8
<< nsubdiff >>
rect 36 432 89 450
rect 36 415 54 432
rect 71 415 89 432
rect 36 397 89 415
<< psubdiffcont >>
rect 54 -8 71 9
<< nsubdiffcont >>
rect 54 415 71 432
<< poly >>
rect 140 400 173 408
rect 140 398 148 400
rect 101 383 148 398
rect 165 383 173 400
rect 101 357 116 383
rect 140 375 173 383
rect 214 400 247 408
rect 214 383 222 400
rect 239 383 247 400
rect 214 375 247 383
rect 214 357 229 375
rect 15 311 48 319
rect 15 294 23 311
rect 40 294 48 311
rect 15 286 48 294
rect 101 287 116 302
rect 24 141 39 286
rect 214 265 229 302
rect 60 250 229 265
rect 60 191 75 250
rect 250 241 265 260
rect 60 176 90 191
rect 216 176 229 191
rect 24 126 90 141
rect 216 126 229 141
rect 250 118 265 199
rect 250 58 265 76
rect 241 50 274 58
rect 241 48 249 50
rect 0 33 249 48
rect 266 48 274 50
rect 266 33 308 48
rect 241 25 274 33
<< polycont >>
rect 148 383 165 400
rect 222 383 239 400
rect 23 294 40 311
rect 249 33 266 50
<< locali >>
rect 0 432 308 445
rect 0 428 54 432
rect 46 415 54 428
rect 71 428 308 432
rect 71 415 90 428
rect 46 407 90 415
rect 73 357 90 407
rect 140 400 173 408
rect 140 383 148 400
rect 165 393 173 400
rect 214 400 247 408
rect 165 383 196 393
rect 140 375 196 383
rect 214 383 222 400
rect 239 383 247 400
rect 214 375 247 383
rect 179 357 196 375
rect 66 349 99 357
rect 66 332 74 349
rect 91 332 99 349
rect 179 349 212 357
rect 66 324 99 332
rect 118 327 151 335
rect 15 311 48 319
rect 15 294 23 311
rect 40 294 48 311
rect 118 310 126 327
rect 143 310 151 327
rect 118 302 151 310
rect 179 332 187 349
rect 204 332 212 349
rect 264 335 281 428
rect 179 324 212 332
rect 231 327 281 335
rect 15 286 48 294
rect 179 241 196 324
rect 231 310 239 327
rect 256 310 281 327
rect 231 302 264 310
rect 90 233 224 241
rect 90 216 98 233
rect 115 216 144 233
rect 161 216 179 233
rect 196 216 224 233
rect 90 208 224 216
rect 266 233 299 241
rect 266 216 274 233
rect 291 216 299 233
rect 266 199 299 216
rect 90 170 204 175
rect 39 167 204 170
rect 39 153 98 167
rect 39 69 56 153
rect 90 150 98 153
rect 115 150 141 167
rect 158 150 179 167
rect 196 150 204 167
rect 90 142 204 150
rect 90 101 245 109
rect 90 84 98 101
rect 115 84 224 101
rect 241 84 245 101
rect 90 76 245 84
rect 267 101 299 117
rect 267 84 275 101
rect 292 84 299 101
rect 267 76 299 84
rect 39 52 71 69
rect 54 17 71 52
rect 241 50 274 58
rect 241 33 249 50
rect 266 33 274 50
rect 241 25 274 33
rect 46 9 79 17
rect 45 -8 54 9
rect 71 -8 80 9
rect 46 -16 79 -8
<< viali >>
rect 54 415 71 432
rect 148 383 165 400
rect 222 383 239 400
rect 23 294 40 311
rect 126 310 143 327
rect 274 216 291 233
rect 98 84 115 101
rect 275 84 292 101
rect 249 33 266 50
rect 54 -8 71 9
<< metal1 >>
rect 45 438 80 441
rect 45 409 48 438
rect 77 409 80 438
rect 45 406 80 409
rect 142 400 171 406
rect 142 391 148 400
rect 56 383 148 391
rect 165 383 171 400
rect 56 377 171 383
rect 216 400 245 406
rect 216 383 222 400
rect 239 383 245 400
rect 216 377 245 383
rect 56 375 143 377
rect 56 319 72 375
rect 15 311 72 319
rect 15 294 23 311
rect 40 294 72 311
rect 120 327 149 333
rect 222 327 239 377
rect 120 310 126 327
rect 143 310 239 327
rect 120 304 149 310
rect 15 286 72 294
rect 126 139 143 304
rect 215 239 250 242
rect 215 210 218 239
rect 247 233 250 239
rect 268 233 297 239
rect 247 216 274 233
rect 291 216 297 233
rect 247 210 250 216
rect 268 210 297 216
rect 215 207 250 210
rect 98 125 143 139
rect 98 107 115 125
rect 136 107 171 110
rect 92 101 121 107
rect 92 84 98 101
rect 115 84 121 101
rect 92 78 121 84
rect 136 78 139 107
rect 168 101 171 107
rect 269 101 298 107
rect 168 84 275 101
rect 292 84 298 101
rect 168 78 171 84
rect 269 78 298 84
rect 136 75 171 78
rect 243 50 272 56
rect 243 48 249 50
rect 0 33 249 48
rect 266 48 272 50
rect 266 33 308 48
rect 243 27 272 33
rect 45 15 80 18
rect 45 -14 48 15
rect 77 -14 80 15
rect 45 -17 80 -14
<< via1 >>
rect 48 432 77 438
rect 48 415 54 432
rect 54 415 71 432
rect 71 415 77 432
rect 48 409 77 415
rect 218 210 247 239
rect 139 78 168 107
rect 48 9 77 15
rect 48 -8 54 9
rect 54 -8 71 9
rect 71 -8 77 9
rect 48 -14 77 -8
<< metal2 >>
rect 40 441 85 446
rect 40 406 45 441
rect 80 406 85 441
rect 40 401 85 406
rect 136 110 150 468
rect 224 242 238 468
rect 215 239 250 242
rect 215 210 218 239
rect 247 210 250 239
rect 215 207 250 210
rect 136 107 171 110
rect 136 78 139 107
rect 168 78 171 107
rect 136 75 171 78
rect 40 18 85 23
rect 40 -17 45 18
rect 80 -17 85 18
rect 40 -22 85 -17
rect 136 -24 150 75
rect 224 -24 238 207
<< via2 >>
rect 45 438 80 441
rect 45 409 48 438
rect 48 409 77 438
rect 77 409 80 438
rect 45 406 80 409
rect 45 15 80 18
rect 45 -14 48 15
rect 48 -14 77 15
rect 77 -14 80 15
rect 45 -17 80 -14
<< metal3 >>
rect 0 441 308 450
rect 0 420 45 441
rect 36 406 45 420
rect 80 420 308 441
rect 80 406 89 420
rect 36 397 89 406
rect 38 18 87 25
rect 38 15 45 18
rect 0 -15 45 15
rect 38 -17 45 -15
rect 80 15 87 18
rect 80 -15 308 15
rect 80 -17 86 -15
rect 38 -24 86 -17
<< labels >>
flabel locali s 186 340 200 353 0 FreeSans 80 0 0 0 Q_bar
flabel locali s 120 312 134 325 0 FreeSans 80 0 0 0 Q
flabel metal2 s 142 84 159 99 0 FreeSans 200 0 0 0 bl
port 1 nsew
flabel metal2 s 222 214 239 229 0 FreeSans 200 0 0 0 br
port 2 nsew
flabel metal1 s 252 36 269 51 0 FreeSans 200 0 0 0 wl
port 3 nsew
flabel metal3 s 55 421 72 436 0 FreeSans 200 0 0 0 vdd
port 4 nsew
flabel metal3 s 51 -9 68 6 0 FreeSans 200 0 0 0 gnd
port 5 nsew
<< properties >>
string FIXED_BBOX 0 0 308 435
<< end >>
