magic
tech sky130A
timestamp 1606124407
<< nwell >>
rect -31 680 637 683
rect -31 550 666 680
rect -31 458 667 550
rect -29 287 667 458
<< nmos >>
rect 30 25 45 67
rect 218 25 233 67
rect 560 -16 575 68
<< pmos >>
rect 30 308 45 434
rect 218 308 233 434
rect 543 308 558 363
<< ndiff >>
rect -10 55 30 67
rect -10 38 -1 55
rect 16 38 30 55
rect -10 25 30 38
rect 45 55 85 67
rect 45 38 59 55
rect 76 38 85 55
rect 45 25 85 38
rect 178 55 218 67
rect 178 38 187 55
rect 204 38 218 55
rect 178 25 218 38
rect 233 55 321 67
rect 233 38 294 55
rect 311 38 321 55
rect 233 25 321 38
rect 488 55 560 68
rect 488 38 497 55
rect 514 38 560 55
rect 488 -16 560 38
rect 575 11 649 68
rect 575 -6 623 11
rect 640 -6 649 11
rect 575 -16 649 -6
<< pdiff >>
rect -10 420 30 434
rect -10 403 -1 420
rect 16 403 30 420
rect -10 308 30 403
rect 45 338 85 434
rect 45 321 59 338
rect 76 321 85 338
rect 45 308 85 321
rect 118 420 218 434
rect 118 403 127 420
rect 144 403 218 420
rect 118 366 218 403
rect 118 349 127 366
rect 144 349 218 366
rect 118 308 218 349
rect 233 371 321 434
rect 233 354 260 371
rect 277 354 294 371
rect 311 354 321 371
rect 233 337 321 354
rect 233 320 260 337
rect 277 320 294 337
rect 311 320 321 337
rect 233 308 321 320
rect 488 337 543 363
rect 488 320 497 337
rect 514 320 543 337
rect 488 308 543 320
rect 558 338 649 363
rect 558 321 623 338
rect 640 321 649 338
rect 558 308 649 321
<< ndiffc >>
rect -1 38 16 55
rect 59 38 76 55
rect 187 38 204 55
rect 294 38 311 55
rect 497 38 514 55
rect 623 -6 640 11
<< pdiffc >>
rect -1 403 16 420
rect 59 321 76 338
rect 127 403 144 420
rect 127 349 144 366
rect 260 354 277 371
rect 294 354 311 371
rect 260 320 277 337
rect 294 320 311 337
rect 497 320 514 337
rect 623 321 640 338
<< psubdiff >>
rect 51 -57 92 -45
rect 51 -74 63 -57
rect 80 -74 92 -57
rect 51 -86 92 -74
<< nsubdiff >>
rect 54 643 107 661
rect 54 626 72 643
rect 89 626 107 643
rect 54 608 107 626
<< psubdiffcont >>
rect 63 -74 80 -57
<< nsubdiffcont >>
rect 72 626 89 643
<< poly >>
rect 30 434 45 451
rect 218 434 233 452
rect 543 363 558 379
rect 30 285 45 308
rect -60 270 45 285
rect -60 103 -45 270
rect 218 155 233 308
rect 543 293 558 308
rect 200 147 233 155
rect 200 130 208 147
rect 225 130 233 147
rect 200 122 233 130
rect -60 88 45 103
rect 30 67 45 88
rect 218 67 233 122
rect 560 68 575 81
rect 30 10 45 25
rect 218 10 233 25
rect 560 -50 575 -16
<< polycont >>
rect 208 130 225 147
<< locali >>
rect 64 650 97 651
rect -9 643 155 650
rect -9 626 72 643
rect 89 626 155 643
rect -9 617 155 626
rect -9 420 24 617
rect 128 428 155 617
rect -9 403 -1 420
rect 16 403 24 420
rect -9 395 24 403
rect 119 420 181 428
rect 119 403 127 420
rect 144 403 181 420
rect 119 366 181 403
rect 119 349 127 366
rect 144 349 181 366
rect 51 338 84 346
rect 119 341 181 349
rect 252 371 319 430
rect 252 354 260 371
rect 277 354 294 371
rect 311 354 319 371
rect 252 341 319 354
rect 489 341 522 346
rect 51 321 59 338
rect 76 321 84 338
rect 51 313 84 321
rect 252 337 522 341
rect 252 320 260 337
rect 277 320 294 337
rect 311 321 497 337
rect 311 320 319 321
rect 60 296 78 313
rect 252 312 319 320
rect 60 276 160 296
rect 140 150 160 276
rect 200 150 233 155
rect 140 147 233 150
rect 140 130 208 147
rect 225 130 233 147
rect 140 105 160 130
rect 200 122 233 130
rect 60 86 160 105
rect 60 63 78 86
rect -9 55 24 63
rect -9 38 -1 55
rect 16 38 24 55
rect -9 30 24 38
rect 51 55 84 63
rect 51 38 59 55
rect 76 38 84 55
rect 51 30 84 38
rect 179 55 212 63
rect 179 38 187 55
rect 204 38 212 55
rect 179 30 212 38
rect 286 60 319 63
rect 400 60 454 321
rect 489 320 497 321
rect 514 320 522 337
rect 489 312 522 320
rect 615 341 648 346
rect 615 338 843 341
rect 615 321 623 338
rect 640 321 843 338
rect 615 313 648 321
rect 489 60 522 63
rect 286 55 522 60
rect 286 38 294 55
rect 311 40 497 55
rect 311 38 319 40
rect 286 30 319 38
rect 489 38 497 40
rect 514 38 522 55
rect 489 30 522 38
rect 0 -57 20 30
rect 55 -57 88 -49
rect 183 -57 203 30
rect 615 11 648 19
rect 823 11 843 321
rect 615 -6 623 11
rect 640 -6 843 11
rect 615 -9 843 -6
rect 615 -14 648 -9
rect -11 -74 63 -57
rect 80 -74 203 -57
rect 55 -82 88 -74
<< viali >>
rect 72 626 89 643
rect 63 -74 80 -57
<< metal1 >>
rect 54 643 107 661
rect 54 626 72 643
rect 89 626 107 643
rect 54 608 107 626
rect 51 -57 92 -45
rect 51 -74 63 -57
rect 80 -74 92 -57
rect 51 -86 92 -74
<< labels >>
flabel poly s 563 12 574 20 0 FreeSans 200 0 0 0 en
port 6 nsew
flabel locali s 823 136 833 149 0 FreeSans 200 0 0 0 out
port 0 nsew
flabel poly s 546 311 552 317 0 FreeSans 200 0 0 0 enb
port 1 nsew
flabel metal1 s 66 -71 75 -63 0 FreeSans 200 0 0 0 gnd
port 2 nsew
flabel locali s 211 133 222 141 0 FreeSans 200 0 0 0 net1
flabel poly s 33 80 42 90 0 FreeSans 200 0 0 0 in
port 4 nsew
flabel locali s 331 325 345 332 0 FreeSans 200 0 0 0 net2
flabel metal1 s 75 629 86 637 0 FreeSans 200 0 0 0 vdd
port 5 nsew
<< end >>
