Sense Amplifier
.lib "../../sky130_fd_pr/models/sky130.lib.spice" tt

XM1 out bl 3 gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42
XM2 2 blb 3 gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42
XM3 out 2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1
XM4 2 2 vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.55
XM5 3 rd_en gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1
XM6 dout out vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.55
XM7 dout out gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42 

V1 vdd gnd dc 1.8v
V2 blb 0 pulse 1.8 0 0 60ps 60ps 1ns 2ns
V3 bl 0 pulse 0 1.8 0 60ps 60ps 1ns 2ns
V4 rd_en 0 pulse 0 1.8 0 60ps 60ps 5ns 10ns

.tran 0.1p 20n
.control
run
plot V(rd_en)+6 V(bl)+4 V(blb)+2 V(dout) 
.endc
.end
