magic
tech sky130A
timestamp 1616272782
<< nwell >>
rect 70 428 517 635
rect 701 428 1294 635
<< nmos >>
rect 138 81 153 123
rect 288 81 303 123
rect 434 81 449 123
rect 598 64 613 148
rect 769 81 784 123
rect 919 81 934 123
rect 1065 81 1080 123
rect 1229 49 1244 133
<< pmos >>
rect 138 448 153 503
rect 288 448 303 503
rect 434 448 449 503
rect 769 448 784 503
rect 919 448 934 503
rect 1065 448 1080 503
<< ndiff >>
rect 88 111 138 123
rect 88 94 103 111
rect 120 94 138 111
rect 88 81 138 94
rect 153 111 203 123
rect 153 94 171 111
rect 188 94 203 111
rect 153 81 203 94
rect 238 111 288 123
rect 238 94 253 111
rect 270 94 288 111
rect 238 81 288 94
rect 303 111 353 123
rect 303 94 321 111
rect 338 94 353 111
rect 303 81 353 94
rect 384 111 434 123
rect 384 94 399 111
rect 416 94 434 111
rect 384 81 434 94
rect 449 111 499 123
rect 449 94 467 111
rect 484 94 499 111
rect 449 81 499 94
rect 548 111 598 148
rect 548 94 563 111
rect 580 94 598 111
rect 548 64 598 94
rect 613 111 663 148
rect 613 94 631 111
rect 648 94 663 111
rect 613 64 663 94
rect 719 111 769 123
rect 719 94 734 111
rect 751 94 769 111
rect 719 81 769 94
rect 784 111 834 123
rect 784 94 802 111
rect 819 94 834 111
rect 784 81 834 94
rect 869 111 919 123
rect 869 94 884 111
rect 901 94 919 111
rect 869 81 919 94
rect 934 111 973 123
rect 934 94 952 111
rect 969 94 973 111
rect 934 81 973 94
rect 1018 111 1065 123
rect 1018 94 1030 111
rect 1047 94 1065 111
rect 1018 81 1065 94
rect 1080 111 1130 123
rect 1080 94 1098 111
rect 1115 94 1130 111
rect 1080 81 1130 94
rect 1179 111 1229 133
rect 1179 94 1194 111
rect 1211 94 1229 111
rect 1179 49 1229 94
rect 1244 111 1294 133
rect 1244 94 1262 111
rect 1279 94 1294 111
rect 1244 49 1294 94
<< pdiff >>
rect 88 484 138 503
rect 88 467 103 484
rect 120 467 138 484
rect 88 448 138 467
rect 153 484 203 503
rect 153 467 171 484
rect 188 467 203 484
rect 153 448 203 467
rect 238 484 288 503
rect 238 467 253 484
rect 270 467 288 484
rect 238 448 288 467
rect 303 484 353 503
rect 303 467 321 484
rect 338 467 353 484
rect 303 448 353 467
rect 384 484 434 503
rect 384 467 399 484
rect 416 467 434 484
rect 384 448 434 467
rect 449 484 499 503
rect 449 467 467 484
rect 484 467 499 484
rect 449 448 499 467
rect 719 484 769 503
rect 719 467 734 484
rect 751 467 769 484
rect 719 448 769 467
rect 784 484 834 503
rect 784 467 802 484
rect 819 467 834 484
rect 784 448 834 467
rect 869 484 919 503
rect 869 467 884 484
rect 901 467 919 484
rect 869 448 919 467
rect 934 484 984 503
rect 934 467 952 484
rect 969 467 984 484
rect 934 448 984 467
rect 1015 484 1065 503
rect 1015 467 1030 484
rect 1047 467 1065 484
rect 1015 448 1065 467
rect 1080 484 1130 503
rect 1080 467 1098 484
rect 1115 467 1130 484
rect 1080 448 1130 467
<< ndiffc >>
rect 103 94 120 111
rect 171 94 188 111
rect 253 94 270 111
rect 321 94 338 111
rect 399 94 416 111
rect 467 94 484 111
rect 563 94 580 111
rect 631 94 648 111
rect 734 94 751 111
rect 802 94 819 111
rect 884 94 901 111
rect 952 94 969 111
rect 1030 94 1047 111
rect 1098 94 1115 111
rect 1194 94 1211 111
rect 1262 94 1279 111
<< pdiffc >>
rect 103 467 120 484
rect 171 467 188 484
rect 253 467 270 484
rect 321 467 338 484
rect 399 467 416 484
rect 467 467 484 484
rect 734 467 751 484
rect 802 467 819 484
rect 884 467 901 484
rect 952 467 969 484
rect 1030 467 1047 484
rect 1098 467 1115 484
<< psubdiff >>
rect 126 8 167 20
rect 126 -9 138 8
rect 155 -9 167 8
rect 126 -21 167 -9
rect 276 8 317 20
rect 276 -9 288 8
rect 305 -9 317 8
rect 276 -21 317 -9
rect 422 8 463 20
rect 422 -9 434 8
rect 451 -9 463 8
rect 422 -21 463 -9
rect 586 8 627 20
rect 586 -9 598 8
rect 615 -9 627 8
rect 586 -21 627 -9
rect 757 8 798 20
rect 757 -9 769 8
rect 786 -9 798 8
rect 757 -21 798 -9
rect 907 8 948 20
rect 907 -9 919 8
rect 936 -9 948 8
rect 907 -21 948 -9
rect 1053 8 1094 20
rect 1053 -9 1065 8
rect 1082 -9 1094 8
rect 1053 -21 1094 -9
rect 1217 8 1258 20
rect 1217 -9 1229 8
rect 1246 -9 1258 8
rect 1217 -21 1258 -9
<< nsubdiff >>
rect 113 590 166 608
rect 113 573 131 590
rect 148 573 166 590
rect 113 555 166 573
rect 263 590 316 608
rect 263 573 281 590
rect 298 573 316 590
rect 263 555 316 573
rect 409 590 462 608
rect 409 573 427 590
rect 444 573 462 590
rect 409 555 462 573
rect 744 590 797 608
rect 744 573 762 590
rect 779 573 797 590
rect 744 555 797 573
rect 894 590 947 608
rect 894 573 912 590
rect 929 573 947 590
rect 894 555 947 573
rect 1040 590 1093 608
rect 1040 573 1058 590
rect 1075 573 1093 590
rect 1040 555 1093 573
rect 1178 590 1231 608
rect 1178 573 1196 590
rect 1213 573 1231 590
rect 1178 555 1231 573
<< psubdiffcont >>
rect 138 -9 155 8
rect 288 -9 305 8
rect 434 -9 451 8
rect 598 -9 615 8
rect 769 -9 786 8
rect 919 -9 936 8
rect 1065 -9 1082 8
rect 1229 -9 1246 8
<< nsubdiffcont >>
rect 131 573 148 590
rect 281 573 298 590
rect 427 573 444 590
rect 762 573 779 590
rect 912 573 929 590
rect 1058 573 1075 590
rect 1196 573 1213 590
<< poly >>
rect 138 503 153 518
rect 288 503 303 518
rect 434 503 449 518
rect 769 503 784 518
rect 919 503 934 518
rect 1065 503 1080 518
rect 80 191 113 199
rect 80 174 88 191
rect 105 189 113 191
rect 138 189 153 448
rect 288 384 303 448
rect 279 376 312 384
rect 279 359 287 376
rect 304 359 312 376
rect 279 351 312 359
rect 105 174 153 189
rect 80 166 113 174
rect 138 123 153 174
rect 288 123 303 351
rect 434 252 449 448
rect 711 375 744 383
rect 711 358 719 375
rect 736 373 744 375
rect 769 373 784 448
rect 919 384 934 448
rect 736 358 784 373
rect 711 350 744 358
rect 416 244 449 252
rect 416 227 424 244
rect 441 227 449 244
rect 416 219 449 227
rect 434 123 449 219
rect 530 191 563 199
rect 530 174 538 191
rect 555 189 563 191
rect 555 174 613 189
rect 530 166 563 174
rect 598 148 613 174
rect 138 66 153 81
rect 288 66 303 81
rect 434 66 449 81
rect 769 123 784 358
rect 910 376 943 384
rect 910 359 918 376
rect 935 359 943 376
rect 910 351 943 359
rect 919 123 934 351
rect 1065 265 1080 448
rect 1047 257 1080 265
rect 1047 240 1055 257
rect 1072 240 1080 257
rect 1047 232 1080 240
rect 1065 123 1080 232
rect 1161 191 1194 199
rect 1161 174 1169 191
rect 1186 189 1194 191
rect 1186 174 1244 189
rect 1161 166 1194 174
rect 1229 133 1244 174
rect 769 66 784 81
rect 919 66 934 81
rect 1065 66 1080 81
rect 598 49 613 64
rect 1229 34 1244 49
<< polycont >>
rect 88 174 105 191
rect 287 359 304 376
rect 719 358 736 375
rect 424 227 441 244
rect 538 174 555 191
rect 918 359 935 376
rect 1055 240 1072 257
rect 1169 174 1186 191
<< locali >>
rect 70 591 1294 603
rect 70 590 563 591
rect 70 573 131 590
rect 148 573 188 590
rect 205 573 281 590
rect 298 573 338 590
rect 355 573 427 590
rect 444 573 484 590
rect 501 574 563 590
rect 580 574 622 591
rect 639 574 670 591
rect 687 590 1294 591
rect 687 574 762 590
rect 501 573 762 574
rect 779 573 819 590
rect 836 573 912 590
rect 929 573 969 590
rect 986 573 1058 590
rect 1075 573 1115 590
rect 1132 573 1196 590
rect 1213 573 1253 590
rect 1270 573 1294 590
rect 70 558 1294 573
rect 103 503 123 558
rect 253 503 273 558
rect 734 503 754 558
rect 884 503 904 558
rect 95 484 128 503
rect 95 467 103 484
rect 120 467 128 484
rect 95 459 128 467
rect 163 484 196 503
rect 163 467 171 484
rect 188 467 196 484
rect 163 459 196 467
rect 245 484 278 503
rect 245 467 253 484
rect 270 467 278 484
rect 245 459 278 467
rect 313 484 424 503
rect 313 467 321 484
rect 338 467 399 484
rect 416 467 424 484
rect 313 459 424 467
rect 459 484 492 503
rect 459 467 467 484
rect 484 467 492 484
rect 459 459 492 467
rect 726 484 759 503
rect 726 467 734 484
rect 751 467 759 484
rect 726 459 759 467
rect 794 484 827 503
rect 794 467 802 484
rect 819 467 827 484
rect 794 459 827 467
rect 876 484 909 503
rect 876 467 884 484
rect 901 467 909 484
rect 876 459 909 467
rect 944 484 1055 503
rect 944 467 952 484
rect 969 467 1030 484
rect 1047 467 1055 484
rect 944 459 1055 467
rect 1090 484 1123 503
rect 1090 467 1098 484
rect 1115 467 1123 484
rect 1090 459 1123 467
rect 168 377 188 459
rect 468 434 488 459
rect 461 428 491 434
rect 461 411 468 428
rect 485 411 491 428
rect 461 405 491 411
rect 279 377 312 384
rect 711 377 744 383
rect 168 376 744 377
rect 168 359 287 376
rect 304 375 744 376
rect 304 359 719 375
rect 168 358 719 359
rect 736 358 744 375
rect 168 357 744 358
rect 0 191 30 196
rect 80 191 113 199
rect 0 189 88 191
rect 0 172 7 189
rect 24 174 88 189
rect 105 174 113 191
rect 24 172 113 174
rect 0 171 113 172
rect 0 166 30 171
rect 80 166 113 171
rect 168 119 188 357
rect 279 351 312 357
rect 711 350 744 357
rect 799 377 819 459
rect 1099 434 1119 459
rect 1092 428 1122 434
rect 1092 411 1099 428
rect 1116 411 1122 428
rect 1092 405 1122 411
rect 910 377 943 384
rect 799 376 943 377
rect 799 359 918 376
rect 935 359 943 376
rect 799 357 943 359
rect 631 328 661 334
rect 631 311 638 328
rect 655 311 661 328
rect 631 305 661 311
rect 586 255 616 261
rect 416 249 449 252
rect 586 249 593 255
rect 230 244 260 249
rect 416 244 593 249
rect 230 242 424 244
rect 230 225 237 242
rect 254 227 424 242
rect 441 238 593 244
rect 610 238 616 255
rect 441 232 616 238
rect 441 227 449 232
rect 254 225 449 227
rect 230 224 449 225
rect 230 219 260 224
rect 416 219 449 224
rect 461 195 491 201
rect 461 194 468 195
rect 328 178 468 194
rect 485 194 491 195
rect 530 194 563 199
rect 485 191 563 194
rect 485 178 538 191
rect 328 174 538 178
rect 555 174 563 191
rect 328 119 348 174
rect 461 172 491 174
rect 468 119 488 172
rect 530 166 563 174
rect 633 119 653 305
rect 799 119 819 357
rect 910 351 943 357
rect 984 329 1014 334
rect 1247 329 1277 334
rect 984 328 1277 329
rect 984 311 991 328
rect 1008 311 1254 328
rect 1271 311 1277 328
rect 984 309 1277 311
rect 984 305 1014 309
rect 1247 305 1277 309
rect 1047 257 1080 265
rect 1047 240 1055 257
rect 1072 240 1080 257
rect 1047 232 1080 240
rect 1092 195 1122 201
rect 1092 194 1099 195
rect 948 178 1099 194
rect 1116 194 1122 195
rect 1161 194 1194 199
rect 1116 191 1194 194
rect 1116 178 1169 191
rect 948 174 1169 178
rect 1186 174 1194 191
rect 948 119 968 174
rect 1092 172 1122 174
rect 1098 119 1118 172
rect 1161 166 1194 174
rect 1263 191 1293 197
rect 1263 174 1270 191
rect 1287 174 1293 191
rect 1263 168 1293 174
rect 1263 119 1283 168
rect 95 111 128 119
rect 95 94 103 111
rect 120 94 128 111
rect 95 81 128 94
rect 163 111 196 119
rect 163 94 171 111
rect 188 94 196 111
rect 163 81 196 94
rect 245 111 278 119
rect 245 94 253 111
rect 270 94 278 111
rect 245 81 278 94
rect 313 111 353 119
rect 313 94 321 111
rect 338 94 353 111
rect 313 81 353 94
rect 384 111 424 119
rect 384 94 399 111
rect 416 94 424 111
rect 384 81 424 94
rect 459 111 492 119
rect 459 94 467 111
rect 484 94 492 111
rect 459 81 492 94
rect 555 111 588 119
rect 555 94 563 111
rect 580 94 588 111
rect 555 81 588 94
rect 623 111 656 119
rect 623 94 631 111
rect 648 94 656 111
rect 623 81 656 94
rect 726 111 759 119
rect 726 94 734 111
rect 751 94 759 111
rect 726 81 759 94
rect 794 111 827 119
rect 794 94 802 111
rect 819 94 827 111
rect 794 81 827 94
rect 876 111 909 119
rect 876 94 884 111
rect 901 94 909 111
rect 876 81 909 94
rect 944 111 973 119
rect 944 94 952 111
rect 969 94 973 111
rect 944 81 973 94
rect 1018 111 1055 119
rect 1018 94 1030 111
rect 1047 94 1055 111
rect 1018 81 1055 94
rect 1090 111 1123 119
rect 1090 94 1098 111
rect 1115 94 1123 111
rect 1090 81 1123 94
rect 1186 111 1219 119
rect 1186 94 1194 111
rect 1211 94 1219 111
rect 1186 81 1219 94
rect 1254 111 1287 119
rect 1254 94 1262 111
rect 1279 94 1287 111
rect 1254 81 1287 94
rect 98 16 118 81
rect 253 16 273 81
rect 393 16 413 81
rect 563 16 583 81
rect 729 16 749 81
rect 884 16 904 81
rect 1023 16 1043 81
rect 1194 16 1214 81
rect 70 8 1294 16
rect 70 -9 103 8
rect 120 -9 138 8
rect 155 -9 181 8
rect 198 -9 253 8
rect 270 -9 288 8
rect 305 -9 331 8
rect 348 -9 399 8
rect 416 -9 434 8
rect 451 -9 477 8
rect 494 -9 563 8
rect 580 -9 598 8
rect 615 -9 641 8
rect 658 -9 734 8
rect 751 -9 769 8
rect 786 -9 812 8
rect 829 -9 884 8
rect 901 -9 919 8
rect 936 -9 962 8
rect 979 -9 1030 8
rect 1047 -9 1065 8
rect 1082 -9 1108 8
rect 1125 -9 1194 8
rect 1211 -9 1229 8
rect 1246 -9 1272 8
rect 1289 -9 1294 8
rect 70 -17 1294 -9
<< viali >>
rect 188 573 205 590
rect 338 573 355 590
rect 484 573 501 590
rect 563 574 580 591
rect 622 574 639 591
rect 670 574 687 591
rect 819 573 836 590
rect 969 573 986 590
rect 1115 573 1132 590
rect 1253 573 1270 590
rect 468 411 485 428
rect 7 172 24 189
rect 88 174 105 191
rect 1099 411 1116 428
rect 638 311 655 328
rect 237 225 254 242
rect 424 227 441 244
rect 593 238 610 255
rect 468 178 485 195
rect 991 311 1008 328
rect 1254 311 1271 328
rect 1055 240 1072 257
rect 1099 178 1116 195
rect 1270 174 1287 191
rect 103 -9 120 8
rect 181 -9 198 8
rect 253 -9 270 8
rect 331 -9 348 8
rect 399 -9 416 8
rect 477 -9 494 8
rect 563 -9 580 8
rect 641 -9 658 8
rect 734 -9 751 8
rect 812 -9 829 8
rect 884 -9 901 8
rect 962 -9 979 8
rect 1030 -9 1047 8
rect 1108 -9 1125 8
rect 1194 -9 1211 8
rect 1272 -9 1289 8
<< metal1 >>
rect 70 591 1294 603
rect 70 590 563 591
rect 70 573 188 590
rect 205 573 338 590
rect 355 573 484 590
rect 501 574 563 590
rect 580 574 622 591
rect 639 574 670 591
rect 687 590 1294 591
rect 687 574 819 590
rect 501 573 819 574
rect 836 573 969 590
rect 986 573 1115 590
rect 1132 573 1253 590
rect 1270 573 1294 590
rect 70 558 1294 573
rect 461 428 491 434
rect 461 411 468 428
rect 485 411 491 428
rect 230 244 260 249
rect 57 242 260 244
rect 57 225 237 242
rect 254 225 260 242
rect 57 224 260 225
rect 230 219 260 224
rect 418 244 447 250
rect 418 227 424 244
rect 441 227 447 244
rect 418 221 447 227
rect 0 189 30 196
rect 0 172 7 189
rect 24 172 30 189
rect 0 166 30 172
rect 82 191 111 197
rect 82 174 88 191
rect 105 174 111 191
rect 82 168 111 174
rect 461 195 491 411
rect 1092 428 1122 434
rect 1092 411 1099 428
rect 1116 411 1122 428
rect 1092 405 1122 411
rect 631 328 1014 334
rect 631 311 638 328
rect 655 311 991 328
rect 1008 311 1014 328
rect 631 305 1014 311
rect 1047 261 1080 265
rect 586 257 1080 261
rect 586 255 1055 257
rect 586 238 593 255
rect 610 240 1055 255
rect 1072 240 1080 257
rect 610 238 1080 240
rect 586 232 1080 238
rect 1096 201 1122 405
rect 1247 328 1277 334
rect 1247 311 1254 328
rect 1271 311 1277 328
rect 1247 305 1277 311
rect 461 178 468 195
rect 485 178 491 195
rect 461 172 491 178
rect 1092 195 1122 201
rect 1092 178 1099 195
rect 1116 178 1122 195
rect 1092 172 1122 178
rect 1263 191 1293 197
rect 1263 174 1270 191
rect 1287 174 1293 191
rect 1263 168 1293 174
rect 70 8 1294 16
rect 70 -9 103 8
rect 120 -9 181 8
rect 198 -9 253 8
rect 270 -9 331 8
rect 348 -9 399 8
rect 416 -9 477 8
rect 494 -9 563 8
rect 580 -9 641 8
rect 658 -9 734 8
rect 751 -9 812 8
rect 829 -9 884 8
rect 901 -9 962 8
rect 979 -9 1030 8
rect 1047 -9 1108 8
rect 1125 -9 1194 8
rect 1211 -9 1272 8
rect 1289 -9 1294 8
rect 70 -17 1294 -9
<< labels >>
flabel locali s 824 363 834 374 0 FreeSans 200 0 0 0 net3
flabel locali s 1102 182 1112 193 0 FreeSans 200 0 0 0 net4
flabel locali s 470 180 480 191 0 FreeSans 200 0 0 0 net2
flabel locali s 359 470 369 481 0 FreeSans 200 0 0 0 net5
flabel locali s 991 470 1001 481 0 FreeSans 200 0 0 0 net6
flabel locali s 176 304 186 315 0 FreeSans 200 0 0 0 net1
flabel metal1 s 10 175 23 187 0 FreeSans 400 0 0 0 din
port 6 nsew
flabel metal1 s 1274 179 1284 188 0 FreeSans 400 0 0 0 bl
port 7 nsew
flabel metal1 s 1257 315 1267 324 0 FreeSans 400 0 0 0 br
port 8 nsew
flabel metal1 s 425 228 438 242 0 FreeSans 400 0 0 0 en
port 9 nsew
flabel metal1 s 505 -12 544 7 0 FreeSans 400 0 0 0 gnd
port 11 nsew
flabel metal1 s 521 571 560 592 0 FreeSans 400 0 0 0 vdd
port 10 nsew
<< properties >>
string FIXED_BBOX 0 0 1294 582
<< end >>
