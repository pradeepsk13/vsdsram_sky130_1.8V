6T SRAM Cell (READ)

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

**********Access Transistors********************
XM1 bl wl q gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42
XM2 blb wl qb gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42


***********Inverter 1*****************************
XM3 q qb vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.55
XM4 q qb gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1.26

*************Inverter 2 ***************************
XM5 qb q vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.55
XM6 qb q gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1.26

V1 vdd gnd dc 1.8v
Vwl wl gnd pulse 0 1.8 0 60ps 60ps 20ns 40ns
Vq q gnd pulse 0 1.8 0 60ps 60ps 5ns 10ns

.tran 0.1n 100n 
.control
run
plot V(wl)+8 V(bl)+2 V(blb) V(q)+6 V(qb)+4
.endc
.end
