magic
tech sky130A
timestamp 1614935929
<< nwell >>
rect 24 188 251 418
<< nmos >>
rect 76 49 91 91
rect 130 49 145 91
rect 174 49 189 91
rect 267 49 282 91
<< pmos >>
rect 76 206 91 332
rect 130 206 145 332
rect 181 206 196 261
<< ndiff >>
rect 51 89 76 91
rect 42 81 76 89
rect 42 64 50 81
rect 67 64 76 81
rect 42 49 76 64
rect 91 81 130 91
rect 91 64 100 81
rect 117 64 130 81
rect 91 49 130 64
rect 145 82 174 91
rect 145 65 151 82
rect 168 65 174 82
rect 145 49 174 65
rect 189 83 267 91
rect 189 66 206 83
rect 223 66 240 83
rect 257 66 267 83
rect 189 49 267 66
rect 282 81 315 91
rect 282 64 290 81
rect 307 64 315 81
rect 282 49 315 64
<< pdiff >>
rect 42 318 76 332
rect 42 301 47 318
rect 64 301 76 318
rect 42 245 76 301
rect 42 228 47 245
rect 64 228 76 245
rect 42 206 76 228
rect 91 312 130 332
rect 91 295 99 312
rect 116 295 130 312
rect 91 245 130 295
rect 91 228 99 245
rect 116 228 130 245
rect 91 206 130 228
rect 145 312 173 332
rect 145 295 151 312
rect 168 295 173 312
rect 145 261 173 295
rect 145 245 181 261
rect 145 228 152 245
rect 169 228 181 245
rect 145 206 181 228
rect 196 245 233 261
rect 196 228 208 245
rect 225 228 233 245
rect 196 206 233 228
<< ndiffc >>
rect 50 64 67 81
rect 100 64 117 81
rect 151 65 168 82
rect 206 66 223 83
rect 240 66 257 83
rect 290 64 307 81
<< pdiffc >>
rect 47 301 64 318
rect 47 228 64 245
rect 99 295 116 312
rect 99 228 116 245
rect 151 295 168 312
rect 152 228 169 245
rect 208 228 225 245
<< psubdiff >>
rect 89 9 130 21
rect 89 -8 101 9
rect 118 -8 130 9
rect 89 -20 130 -8
<< nsubdiff >>
rect 43 388 84 400
rect 43 371 55 388
rect 72 371 84 388
rect 43 359 84 371
<< psubdiffcont >>
rect 101 -8 118 9
<< nsubdiffcont >>
rect 55 371 72 388
<< poly >>
rect 76 332 91 346
rect 130 332 145 346
rect 243 306 276 314
rect 243 304 251 306
rect 181 289 251 304
rect 268 304 276 306
rect 268 289 282 304
rect 181 261 196 289
rect 243 281 282 289
rect 6 133 39 139
rect 76 133 91 206
rect 130 188 145 206
rect 181 193 196 206
rect 112 180 145 188
rect 112 163 120 180
rect 137 163 145 180
rect 112 155 145 163
rect 6 131 91 133
rect 6 114 14 131
rect 31 118 91 131
rect 31 114 39 118
rect 6 106 39 114
rect 76 91 91 118
rect 130 91 145 155
rect 166 161 199 169
rect 166 144 174 161
rect 191 144 199 161
rect 166 136 199 144
rect 174 91 189 136
rect 267 91 282 281
rect 76 36 91 49
rect 130 36 145 49
rect 174 36 189 49
rect 267 36 282 49
<< polycont >>
rect 251 289 268 306
rect 120 163 137 180
rect 14 114 31 131
rect 174 144 191 161
<< locali >>
rect 47 388 80 396
rect 0 371 55 388
rect 72 371 124 388
rect 141 371 200 388
rect 217 371 280 388
rect 297 371 320 388
rect 47 363 80 371
rect 42 318 73 332
rect 100 322 117 371
rect 42 301 47 318
rect 64 301 73 318
rect 42 245 73 301
rect 42 228 47 245
rect 64 228 73 245
rect 42 206 73 228
rect 91 312 124 322
rect 91 295 99 312
rect 116 295 124 312
rect 91 245 124 295
rect 91 228 99 245
rect 116 228 124 245
rect 91 206 124 228
rect 145 312 173 322
rect 145 295 151 312
rect 168 295 173 312
rect 145 261 173 295
rect 243 306 276 314
rect 243 289 251 306
rect 268 289 276 306
rect 243 281 276 289
rect 145 245 178 261
rect 145 228 152 245
rect 169 228 178 245
rect 145 206 178 228
rect 200 245 233 261
rect 200 228 208 245
rect 225 228 233 245
rect 200 206 233 228
rect 56 180 73 206
rect 216 196 233 206
rect 112 180 145 188
rect 56 163 120 180
rect 137 163 145 180
rect 216 179 275 196
rect 6 131 39 139
rect 6 114 14 131
rect 31 114 39 131
rect 6 106 39 114
rect 56 89 73 163
rect 112 155 145 163
rect 166 161 199 169
rect 166 144 174 161
rect 191 144 199 161
rect 166 136 199 144
rect 216 91 233 179
rect 42 81 75 89
rect 42 64 50 81
rect 67 64 75 81
rect 42 49 75 64
rect 92 81 125 91
rect 92 64 100 81
rect 117 64 125 81
rect 92 56 125 64
rect 145 82 176 91
rect 145 65 151 82
rect 168 65 176 82
rect 100 17 117 56
rect 145 55 176 65
rect 198 89 248 91
rect 198 83 265 89
rect 198 66 206 83
rect 223 66 240 83
rect 257 66 265 83
rect 198 55 265 66
rect 282 81 315 91
rect 282 64 290 81
rect 307 64 315 81
rect 282 56 315 64
rect 93 9 126 17
rect 298 9 315 56
rect 0 -8 20 9
rect 37 -8 101 9
rect 118 -8 203 9
rect 220 -8 298 9
rect 315 -8 320 9
rect 93 -16 126 -8
<< viali >>
rect 55 371 72 388
rect 124 371 141 388
rect 200 371 217 388
rect 280 371 297 388
rect 251 289 268 306
rect 275 179 292 196
rect 14 114 31 131
rect 174 144 191 161
rect 20 -8 37 9
rect 101 -8 118 9
rect 203 -8 220 9
rect 298 -8 315 9
<< metal1 >>
rect 0 388 320 394
rect 0 371 55 388
rect 72 371 124 388
rect 141 371 200 388
rect 217 371 280 388
rect 297 371 320 388
rect 0 365 320 371
rect 243 311 276 314
rect 243 285 246 311
rect 272 285 276 311
rect 243 281 276 285
rect 0 217 320 232
rect 275 202 290 217
rect 269 196 298 202
rect 269 179 275 196
rect 292 179 298 196
rect 269 173 298 179
rect 166 166 199 169
rect 166 140 169 166
rect 195 140 199 166
rect 8 131 37 137
rect 166 136 199 140
rect 8 120 14 131
rect 0 114 14 120
rect 31 120 37 131
rect 31 114 320 120
rect 0 106 320 114
rect 0 9 320 15
rect 0 -8 20 9
rect 37 -8 101 9
rect 118 -8 203 9
rect 220 -8 298 9
rect 315 -8 320 9
rect 0 -14 320 -8
<< via1 >>
rect 246 306 272 311
rect 246 289 251 306
rect 251 289 268 306
rect 268 289 272 306
rect 246 285 272 289
rect 169 161 195 166
rect 169 144 174 161
rect 174 144 191 161
rect 191 144 195 161
rect 169 140 195 144
<< metal2 >>
rect 166 169 180 418
rect 243 314 257 418
rect 243 311 276 314
rect 243 285 246 311
rect 272 285 276 311
rect 243 281 276 285
rect 166 166 199 169
rect 166 140 169 166
rect 195 140 199 166
rect 166 136 199 140
rect 166 -22 180 136
rect 243 -22 257 281
<< labels >>
flabel metal1 s 56 373 69 385 0 FreeSans 200 0 0 0 vdd
port 0 nsew
flabel metal1 s 102 -6 115 6 0 FreeSans 200 0 0 0 gnd
port 2 nsew
flabel metal1 s 278 183 288 192 0 FreeSans 200 0 0 0 out
port 6 nsew
flabel metal2 s 177 149 187 158 0 FreeSans 200 0 0 0 en
port 8 nsew
flabel metal2 s 254 294 264 303 0 FreeSans 200 0 0 0 enb
port 10 nsew
flabel metal1 s 15 115 29 128 0 FreeSans 200 0 0 0 in
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 320 380
<< end >>
