magic
tech sky130A
timestamp 1617114508
<< nwell >>
rect 0 294 308 555
<< nmos >>
rect 52 610 67 652
rect 102 610 117 652
rect 226 611 241 653
rect 52 216 67 258
rect 102 216 117 258
rect 226 196 241 238
rect 71 50 86 134
rect 226 48 241 132
<< pmos >>
rect 52 480 67 535
rect 102 480 117 535
rect 226 480 241 535
rect 52 314 67 369
rect 102 314 117 369
rect 226 314 241 369
<< ndiff >>
rect 18 639 52 652
rect 18 622 26 639
rect 43 622 52 639
rect 18 610 52 622
rect 67 639 102 652
rect 67 622 76 639
rect 93 622 102 639
rect 67 610 102 622
rect 117 639 151 652
rect 117 622 126 639
rect 143 622 151 639
rect 117 610 151 622
rect 192 640 226 653
rect 192 623 200 640
rect 217 623 226 640
rect 192 611 226 623
rect 241 640 275 653
rect 241 623 250 640
rect 267 623 275 640
rect 241 611 275 623
rect 18 246 52 258
rect 18 229 26 246
rect 43 229 52 246
rect 18 216 52 229
rect 67 246 102 258
rect 67 229 76 246
rect 93 229 102 246
rect 67 216 102 229
rect 117 246 151 258
rect 117 229 126 246
rect 143 229 151 246
rect 117 216 151 229
rect 192 226 226 238
rect 192 209 200 226
rect 217 209 226 226
rect 192 196 226 209
rect 241 226 275 238
rect 241 209 250 226
rect 267 209 275 226
rect 241 196 275 209
rect 21 118 71 134
rect 21 101 37 118
rect 54 101 71 118
rect 21 75 71 101
rect 21 58 37 75
rect 54 58 71 75
rect 21 50 71 58
rect 86 123 136 134
rect 86 106 111 123
rect 128 106 136 123
rect 86 78 136 106
rect 86 61 111 78
rect 128 61 136 78
rect 86 50 136 61
rect 176 119 226 132
rect 176 102 195 119
rect 212 102 226 119
rect 176 81 226 102
rect 176 64 195 81
rect 212 64 226 81
rect 176 48 226 64
rect 241 73 291 132
rect 241 56 258 73
rect 275 56 291 73
rect 241 48 291 56
<< pdiff >>
rect 18 516 52 535
rect 18 499 29 516
rect 46 499 52 516
rect 18 480 52 499
rect 67 516 102 535
rect 67 499 76 516
rect 93 499 102 516
rect 67 480 102 499
rect 117 516 151 535
rect 117 499 126 516
rect 143 499 151 516
rect 117 480 151 499
rect 192 516 226 535
rect 192 499 200 516
rect 217 499 226 516
rect 192 480 226 499
rect 241 516 275 535
rect 241 499 250 516
rect 267 499 275 516
rect 241 480 275 499
rect 18 350 52 369
rect 18 333 26 350
rect 43 333 52 350
rect 18 314 52 333
rect 67 350 102 369
rect 67 333 76 350
rect 93 333 102 350
rect 67 314 102 333
rect 117 350 151 369
rect 117 333 126 350
rect 143 333 151 350
rect 117 314 151 333
rect 192 350 226 369
rect 192 333 200 350
rect 217 333 226 350
rect 192 314 226 333
rect 241 350 275 369
rect 241 333 250 350
rect 267 333 275 350
rect 241 314 275 333
<< ndiffc >>
rect 26 622 43 639
rect 76 622 93 639
rect 126 622 143 639
rect 200 623 217 640
rect 250 623 267 640
rect 26 229 43 246
rect 76 229 93 246
rect 126 229 143 246
rect 200 209 217 226
rect 250 209 267 226
rect 37 101 54 118
rect 37 58 54 75
rect 111 106 128 123
rect 111 61 128 78
rect 195 102 212 119
rect 195 64 212 81
rect 258 56 275 73
<< pdiffc >>
rect 29 499 46 516
rect 76 499 93 516
rect 126 499 143 516
rect 200 499 217 516
rect 250 499 267 516
rect 26 333 43 350
rect 76 333 93 350
rect 126 333 143 350
rect 200 333 217 350
rect 250 333 267 350
<< psubdiff >>
rect 63 716 104 728
rect 63 699 75 716
rect 92 699 104 716
rect 63 687 104 699
rect 172 716 213 728
rect 172 699 184 716
rect 201 699 213 716
rect 172 687 213 699
rect 180 9 221 21
rect 180 -8 192 9
rect 209 -8 221 9
rect 180 -20 221 -8
<< nsubdiff >>
rect 188 437 229 449
rect 188 420 200 437
rect 217 420 229 437
rect 188 408 229 420
<< psubdiffcont >>
rect 75 699 92 716
rect 184 699 201 716
rect 192 -8 209 9
<< nsubdiffcont >>
rect 200 420 217 437
<< poly >>
rect 52 652 67 667
rect 102 652 117 667
rect 226 653 241 668
rect 52 591 67 610
rect 34 583 67 591
rect 34 566 42 583
rect 59 566 67 583
rect 34 558 67 566
rect 52 535 67 558
rect 102 575 117 610
rect 172 577 205 585
rect 172 575 180 577
rect 102 560 180 575
rect 197 560 205 577
rect 102 535 117 560
rect 172 552 205 560
rect 226 535 241 611
rect 52 369 67 480
rect 102 465 117 480
rect 226 471 241 480
rect 140 455 241 471
rect 140 408 155 455
rect 102 392 155 408
rect 102 369 117 392
rect 226 369 241 384
rect 52 258 67 314
rect 102 289 117 314
rect 172 289 205 297
rect 102 274 180 289
rect 102 258 117 274
rect 172 272 180 274
rect 197 272 205 289
rect 172 264 205 272
rect 226 292 241 314
rect 226 284 259 292
rect 226 267 234 284
rect 251 267 259 284
rect 226 259 259 267
rect 226 238 241 259
rect 52 201 67 216
rect 102 201 117 216
rect 226 181 241 196
rect 16 171 49 179
rect 16 154 24 171
rect 41 154 86 171
rect 16 146 49 154
rect 71 134 86 154
rect 171 170 204 178
rect 171 153 179 170
rect 196 160 204 170
rect 196 153 241 160
rect 171 145 241 153
rect 226 132 241 145
rect 71 35 86 50
rect 226 33 241 48
<< polycont >>
rect 42 566 59 583
rect 180 560 197 577
rect 180 272 197 289
rect 234 267 251 284
rect 24 154 41 171
rect 179 153 196 170
<< locali >>
rect 67 716 100 724
rect 67 699 75 716
rect 92 699 100 716
rect 67 691 100 699
rect 176 716 209 724
rect 176 699 184 716
rect 201 699 209 716
rect 176 691 209 699
rect 75 647 92 691
rect 186 690 203 691
rect 18 639 51 647
rect 18 622 26 639
rect 43 622 51 639
rect 18 614 51 622
rect 68 639 101 647
rect 68 622 76 639
rect 93 622 101 639
rect 68 614 101 622
rect 118 639 151 647
rect 118 622 126 639
rect 143 622 151 639
rect 118 614 151 622
rect 192 640 225 648
rect 192 623 200 640
rect 217 623 225 640
rect 192 615 225 623
rect 242 640 275 648
rect 242 623 250 640
rect 267 623 275 640
rect 242 615 275 623
rect 34 583 67 591
rect 192 585 209 615
rect 34 566 42 583
rect 59 566 67 583
rect 34 558 67 566
rect 172 577 209 585
rect 172 560 180 577
rect 197 560 209 577
rect 172 552 209 560
rect 18 524 35 535
rect 192 524 209 552
rect 18 516 51 524
rect 18 499 29 516
rect 46 499 51 516
rect 18 480 51 499
rect 68 516 101 524
rect 68 499 76 516
rect 93 499 101 516
rect 68 490 101 499
rect 118 516 151 524
rect 118 499 126 516
rect 143 499 151 516
rect 118 490 151 499
rect 192 516 225 524
rect 192 499 200 516
rect 217 499 225 516
rect 192 489 225 499
rect 242 516 275 524
rect 242 499 250 516
rect 267 499 275 516
rect 242 489 275 499
rect 192 437 225 445
rect 192 420 200 437
rect 217 420 225 437
rect 192 412 225 420
rect 208 411 225 412
rect 257 360 275 489
rect 18 350 51 359
rect 18 333 26 350
rect 43 333 51 350
rect 18 325 51 333
rect 68 350 101 359
rect 68 333 76 350
rect 93 333 101 350
rect 68 325 101 333
rect 118 350 151 359
rect 118 333 126 350
rect 143 333 151 350
rect 118 325 151 333
rect 192 350 225 360
rect 192 333 200 350
rect 217 333 225 350
rect 192 325 225 333
rect 242 350 275 360
rect 242 333 250 350
rect 267 333 275 350
rect 242 325 275 333
rect 18 254 35 325
rect 192 297 209 325
rect 172 289 209 297
rect 172 272 180 289
rect 197 272 209 289
rect 172 264 209 272
rect 18 246 51 254
rect 18 229 26 246
rect 43 229 51 246
rect 18 221 51 229
rect 68 246 101 254
rect 68 229 76 246
rect 93 229 101 246
rect 68 221 101 229
rect 118 246 151 254
rect 118 229 126 246
rect 143 229 151 246
rect 118 221 151 229
rect 192 234 209 264
rect 226 284 259 292
rect 226 267 234 284
rect 251 267 259 284
rect 226 259 259 267
rect 192 226 225 234
rect 16 171 49 179
rect 16 154 24 171
rect 41 154 49 171
rect 16 146 49 154
rect 68 126 86 221
rect 192 209 200 226
rect 217 209 225 226
rect 192 201 225 209
rect 242 226 275 234
rect 242 209 250 226
rect 267 209 275 226
rect 242 201 275 209
rect 171 170 204 178
rect 171 153 179 170
rect 196 153 204 170
rect 171 145 204 153
rect 29 118 86 126
rect 29 101 37 118
rect 54 109 86 118
rect 103 123 136 131
rect 54 101 62 109
rect 29 75 62 101
rect 29 58 37 75
rect 54 58 62 75
rect 29 50 62 58
rect 103 106 111 123
rect 128 106 136 123
rect 103 78 136 106
rect 103 61 111 78
rect 128 61 136 78
rect 103 53 136 61
rect 187 119 220 127
rect 187 102 195 119
rect 212 102 220 119
rect 187 81 220 102
rect 187 64 195 81
rect 212 64 220 81
rect 258 80 275 201
rect 187 56 220 64
rect 250 73 283 80
rect 250 56 258 73
rect 275 56 283 73
rect 250 48 283 56
rect 184 9 217 17
rect 184 -8 192 9
rect 209 -8 217 9
rect 184 -16 217 -8
<< viali >>
rect 75 699 92 716
rect 184 699 201 716
rect 26 622 43 639
rect 126 622 143 639
rect 250 623 267 640
rect 42 566 59 583
rect 126 499 143 516
rect 200 420 217 437
rect 126 333 143 350
rect 26 229 43 246
rect 126 229 143 246
rect 234 267 251 284
rect 24 154 41 171
rect 179 153 196 170
rect 37 101 54 118
rect 37 58 54 75
rect 111 106 128 123
rect 111 61 128 78
rect 195 102 212 119
rect 195 64 212 81
rect 258 56 275 73
rect 192 -8 209 9
<< metal1 >>
rect 175 722 210 725
rect 69 716 98 722
rect 175 716 178 722
rect 207 716 210 722
rect 69 715 75 716
rect 0 699 75 715
rect 92 699 178 716
rect 207 699 308 716
rect 69 693 98 699
rect 175 693 178 699
rect 207 693 210 699
rect 175 690 210 693
rect 16 680 51 683
rect 16 651 19 680
rect 48 651 51 680
rect 16 648 51 651
rect 18 639 51 648
rect 250 646 267 699
rect 120 639 149 645
rect 18 622 26 639
rect 43 622 126 639
rect 143 622 149 639
rect 18 614 51 622
rect 120 616 149 622
rect 244 640 273 646
rect 244 623 250 640
rect 267 623 273 640
rect 244 617 273 623
rect 36 583 65 589
rect 0 566 42 583
rect 59 566 308 583
rect 36 560 65 566
rect 120 516 149 522
rect 120 499 126 516
rect 143 499 149 516
rect 120 493 149 499
rect 125 437 140 493
rect 191 443 226 446
rect 191 437 194 443
rect 223 437 226 443
rect 0 420 194 437
rect 223 420 308 437
rect 125 356 140 420
rect 191 414 194 420
rect 223 414 226 420
rect 191 411 226 414
rect 120 350 149 356
rect 120 333 126 350
rect 143 333 149 350
rect 120 327 149 333
rect 226 284 259 292
rect 0 267 234 284
rect 251 267 308 284
rect 226 259 259 267
rect 20 246 49 252
rect 120 246 149 252
rect 20 229 26 246
rect 43 229 126 246
rect 143 229 149 246
rect 20 223 49 229
rect 120 223 149 229
rect 135 208 200 223
rect 15 177 50 180
rect 15 148 18 177
rect 47 148 50 177
rect 15 145 50 148
rect 88 177 136 180
rect 88 148 91 177
rect 120 148 136 177
rect 185 176 200 208
rect 88 145 136 148
rect 173 170 202 176
rect 173 153 179 170
rect 196 153 202 170
rect 173 147 202 153
rect 31 118 60 124
rect 31 101 37 118
rect 54 101 60 118
rect 31 75 60 101
rect 31 58 37 75
rect 54 58 60 75
rect 31 52 60 58
rect 103 123 136 145
rect 252 128 287 131
rect 252 127 255 128
rect 103 106 111 123
rect 128 106 136 123
rect 103 78 136 106
rect 103 61 111 78
rect 128 61 136 78
rect 103 53 136 61
rect 187 119 255 127
rect 187 102 195 119
rect 212 107 255 119
rect 212 102 220 107
rect 187 81 220 102
rect 252 99 255 107
rect 284 99 287 128
rect 252 96 287 99
rect 187 64 195 81
rect 212 64 220 81
rect 187 56 220 64
rect 252 73 281 79
rect 252 56 258 73
rect 275 56 281 73
rect 37 9 54 52
rect 252 50 281 56
rect 183 15 218 18
rect 183 9 186 15
rect 215 9 218 15
rect 258 9 275 50
rect 0 -8 186 9
rect 215 -8 308 9
rect 183 -14 186 -8
rect 215 -14 218 -8
rect 183 -17 218 -14
<< via1 >>
rect 178 716 207 722
rect 178 699 184 716
rect 184 699 201 716
rect 201 699 207 716
rect 178 693 207 699
rect 19 651 48 680
rect 194 437 223 443
rect 194 420 200 437
rect 200 420 217 437
rect 217 420 223 437
rect 194 414 223 420
rect 18 171 47 177
rect 18 154 24 171
rect 24 154 41 171
rect 41 154 47 171
rect 18 148 47 154
rect 91 148 120 177
rect 255 99 284 128
rect 186 9 215 15
rect 186 -8 192 9
rect 192 -8 209 9
rect 209 -8 215 9
rect 186 -14 215 -8
<< metal2 >>
rect 16 680 51 683
rect 16 651 19 680
rect 48 651 51 680
rect 16 648 51 651
rect 28 180 43 648
rect 88 180 116 733
rect 170 725 215 730
rect 170 690 175 725
rect 210 690 215 725
rect 170 685 215 690
rect 186 446 231 451
rect 186 411 191 446
rect 226 411 231 446
rect 186 406 231 411
rect 14 177 50 180
rect 14 148 18 177
rect 47 148 50 177
rect 14 145 50 148
rect 88 177 123 180
rect 88 148 91 177
rect 120 148 123 177
rect 88 145 123 148
rect 88 -25 116 145
rect 252 131 280 733
rect 252 128 287 131
rect 252 99 255 128
rect 284 99 287 128
rect 252 96 287 99
rect 178 18 223 23
rect 178 -17 183 18
rect 218 -17 223 18
rect 178 -22 223 -17
rect 252 -25 280 96
<< via2 >>
rect 175 722 210 725
rect 175 693 178 722
rect 178 693 207 722
rect 207 693 210 722
rect 175 690 210 693
rect 191 443 226 446
rect 191 414 194 443
rect 194 414 223 443
rect 223 414 226 443
rect 191 411 226 414
rect 183 15 218 18
rect 183 -14 186 15
rect 186 -14 215 15
rect 215 -14 218 15
rect 183 -17 218 -14
<< metal3 >>
rect 168 725 217 733
rect 0 690 175 725
rect 210 690 308 725
rect 168 684 217 690
rect 186 446 231 451
rect 0 411 191 446
rect 226 411 308 446
rect 186 406 231 411
rect 175 18 226 26
rect 0 -17 183 18
rect 218 -17 308 18
rect 175 -25 226 -17
<< labels >>
flabel metal1 s 234 269 251 282 0 FreeSans 200 180 0 0 din
port 0 nsew
flabel metal1 s 50 567 66 581 0 FreeSans 200 0 0 0 en
port 3 nsew
flabel metal2 s 96 156 118 174 0 FreeSans 200 0 0 0 bl
port 1 nsew
flabel metal2 s 256 103 278 121 0 FreeSans 200 0 0 0 br
port 2 nsew
flabel metal3 s 192 -9 213 7 0 FreeSans 200 180 0 0 gnd
port 5 nsew
flabel metal3 s 197 422 214 434 0 FreeSans 200 0 0 0 vdd
port 4 nsew
flabel metal3 s 184 703 205 719 0 FreeSans 200 180 0 0 gnd
<< properties >>
string FIXED_BBOX 0 0 308 708
<< end >>
