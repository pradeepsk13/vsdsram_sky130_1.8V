N-curve Write

.lib "sky130_fd_pr/models/sky130.lib.spice" tt


******Access transistors**********
XM1 gnd wl Q gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42
XM2 blb wl Qb gnd sky130_fd_pr__nfet_01v8 L=0.15 W=0.42

********Cross inverters ********

XM3 Q Qb gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1.26
XM4 Qb Q gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1.26
XM5 Q Qb vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.55
XM6 Qb Q vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.55

V1 vdd gnd dc 1.8V
Vin Q gnd dc 1.8V
Vwl wl gnd dc 1.8v

Vblb blb gnd dc 1.8v

.dc Vin 0 1.8 0.01
.control
run
plot -I(Vin)
.endc
.end
