VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_2_16_sky130A
   CLASS BLOCK ;
   SIZE 65.04 BY 121.62 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  12.04 -11.74 12.56 -11.22 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  25.16 -11.74 25.68 -11.22 ;
      END
   END din0[1]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -14.2 121.1 -13.68 121.62 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -11.74 121.1 -11.22 121.62 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -12.56 121.1 -12.04 121.62 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -13.38 121.1 -12.86 121.62 ;
      END
   END addr0[3]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  -56.84 -9.28 -56.32 -8.76 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER m3 ;
         RECT  -56.84 -6.0 -56.32 -5.48 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER m4 ;
         RECT  -24.86 -11.74 -24.34 -11.22 ;
      END
   END clk0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  64.52 13.68 65.04 14.2 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER m3 ;
         RECT  64.52 10.4 65.04 10.92 ;
      END
   END dout0[1]
   PIN vdd
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -56.02 -7.64 -54.68 -6.3 ;
      END
   END vdd
   PIN gnd
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER m3 ;
         RECT  -56.02 -11.74 -54.68 -10.4 ;
      END
   END gnd
   OBS
   LAYER  m1 ;
      RECT  50.49 33.82 50.84 34.17 ;
      RECT  48.65 33.33 51.25 33.62 ;
      RECT  49.16 33.82 49.51 34.17 ;
      RECT  48.85 34.48 49.14 34.64 ;
      RECT  49.99 36.99 50.28 37.28 ;
      RECT  48.65 38.45 51.25 38.74 ;
      RECT  49.57 36.45 49.86 36.74 ;
      RECT  48.83 34.33 49.16 34.48 ;
      RECT  50.49 43.38 50.84 43.03 ;
      RECT  48.65 43.87 51.25 43.58 ;
      RECT  49.16 43.38 49.51 43.03 ;
      RECT  48.85 42.72 49.14 42.56 ;
      RECT  49.99 40.21 50.28 39.92 ;
      RECT  48.65 38.75 51.25 38.46 ;
      RECT  49.57 40.75 49.86 40.46 ;
      RECT  48.83 42.87 49.16 42.72 ;
      RECT  50.49 44.08 50.84 44.43 ;
      RECT  48.65 43.59 51.25 43.88 ;
      RECT  49.16 44.08 49.51 44.43 ;
      RECT  48.85 44.74 49.14 44.9 ;
      RECT  49.99 47.25 50.28 47.54 ;
      RECT  48.65 48.71 51.25 49.0 ;
      RECT  49.57 46.71 49.86 47.0 ;
      RECT  48.83 44.59 49.16 44.74 ;
      RECT  50.49 53.64 50.84 53.29 ;
      RECT  48.65 54.13 51.25 53.84 ;
      RECT  49.16 53.64 49.51 53.29 ;
      RECT  48.85 52.98 49.14 52.82 ;
      RECT  49.99 50.47 50.28 50.18 ;
      RECT  48.65 49.01 51.25 48.72 ;
      RECT  49.57 51.01 49.86 50.72 ;
      RECT  48.83 53.13 49.16 52.98 ;
      RECT  50.49 54.34 50.84 54.69 ;
      RECT  48.65 53.85 51.25 54.14 ;
      RECT  49.16 54.34 49.51 54.69 ;
      RECT  48.85 55.0 49.14 55.16 ;
      RECT  49.99 57.51 50.28 57.8 ;
      RECT  48.65 58.97 51.25 59.26 ;
      RECT  49.57 56.97 49.86 57.26 ;
      RECT  48.83 54.85 49.16 55.0 ;
      RECT  50.49 63.9 50.84 63.55 ;
      RECT  48.65 64.39 51.25 64.1 ;
      RECT  49.16 63.9 49.51 63.55 ;
      RECT  48.85 63.24 49.14 63.08 ;
      RECT  49.99 60.73 50.28 60.44 ;
      RECT  48.65 59.27 51.25 58.98 ;
      RECT  49.57 61.27 49.86 60.98 ;
      RECT  48.83 63.39 49.16 63.24 ;
      RECT  50.49 64.6 50.84 64.95 ;
      RECT  48.65 64.11 51.25 64.4 ;
      RECT  49.16 64.6 49.51 64.95 ;
      RECT  48.85 65.26 49.14 65.42 ;
      RECT  49.99 67.77 50.28 68.06 ;
      RECT  48.65 69.23 51.25 69.52 ;
      RECT  49.57 67.23 49.86 67.52 ;
      RECT  48.83 65.11 49.16 65.26 ;
      RECT  50.49 74.16 50.84 73.81 ;
      RECT  48.65 74.65 51.25 74.36 ;
      RECT  49.16 74.16 49.51 73.81 ;
      RECT  48.85 73.5 49.14 73.34 ;
      RECT  49.99 70.99 50.28 70.7 ;
      RECT  48.65 69.53 51.25 69.24 ;
      RECT  49.57 71.53 49.86 71.24 ;
      RECT  48.83 73.65 49.16 73.5 ;
      RECT  50.49 74.86 50.84 75.21 ;
      RECT  48.65 74.37 51.25 74.66 ;
      RECT  49.16 74.86 49.51 75.21 ;
      RECT  48.85 75.52 49.14 75.68 ;
      RECT  49.99 78.03 50.28 78.32 ;
      RECT  48.65 79.49 51.25 79.78 ;
      RECT  49.57 77.49 49.86 77.78 ;
      RECT  48.83 75.37 49.16 75.52 ;
      RECT  50.49 84.42 50.84 84.07 ;
      RECT  48.65 84.91 51.25 84.62 ;
      RECT  49.16 84.42 49.51 84.07 ;
      RECT  48.85 83.76 49.14 83.6 ;
      RECT  49.99 81.25 50.28 80.96 ;
      RECT  48.65 79.79 51.25 79.5 ;
      RECT  49.57 81.79 49.86 81.5 ;
      RECT  48.83 83.91 49.16 83.76 ;
      RECT  50.49 85.12 50.84 85.47 ;
      RECT  48.65 84.63 51.25 84.92 ;
      RECT  49.16 85.12 49.51 85.47 ;
      RECT  48.85 85.78 49.14 85.94 ;
      RECT  49.99 88.29 50.28 88.58 ;
      RECT  48.65 89.75 51.25 90.04 ;
      RECT  49.57 87.75 49.86 88.04 ;
      RECT  48.83 85.63 49.16 85.78 ;
      RECT  50.49 94.68 50.84 94.33 ;
      RECT  48.65 95.17 51.25 94.88 ;
      RECT  49.16 94.68 49.51 94.33 ;
      RECT  48.85 94.02 49.14 93.86 ;
      RECT  49.99 91.51 50.28 91.22 ;
      RECT  48.65 90.05 51.25 89.76 ;
      RECT  49.57 92.05 49.86 91.76 ;
      RECT  48.83 94.17 49.16 94.02 ;
      RECT  50.49 95.38 50.84 95.73 ;
      RECT  48.65 94.89 51.25 95.18 ;
      RECT  49.16 95.38 49.51 95.73 ;
      RECT  48.85 96.04 49.14 96.2 ;
      RECT  49.99 98.55 50.28 98.84 ;
      RECT  48.65 100.01 51.25 100.3 ;
      RECT  49.57 98.01 49.86 98.3 ;
      RECT  48.83 95.89 49.16 96.04 ;
      RECT  50.49 104.94 50.84 104.59 ;
      RECT  48.65 105.43 51.25 105.14 ;
      RECT  49.16 104.94 49.51 104.59 ;
      RECT  48.85 104.28 49.14 104.12 ;
      RECT  49.99 101.77 50.28 101.48 ;
      RECT  48.65 100.31 51.25 100.02 ;
      RECT  49.57 102.31 49.86 102.02 ;
      RECT  48.83 104.43 49.16 104.28 ;
      RECT  50.49 105.64 50.84 105.99 ;
      RECT  48.65 105.15 51.25 105.44 ;
      RECT  49.16 105.64 49.51 105.99 ;
      RECT  48.85 106.3 49.14 106.46 ;
      RECT  49.99 108.81 50.28 109.1 ;
      RECT  48.65 110.27 51.25 110.56 ;
      RECT  49.57 108.27 49.86 108.56 ;
      RECT  48.83 106.15 49.16 106.3 ;
      RECT  50.49 115.2 50.84 114.85 ;
      RECT  48.65 115.69 51.25 115.4 ;
      RECT  49.16 115.2 49.51 114.85 ;
      RECT  48.85 114.54 49.14 114.38 ;
      RECT  49.99 112.03 50.28 111.74 ;
      RECT  48.65 110.57 51.25 110.28 ;
      RECT  49.57 112.57 49.86 112.28 ;
      RECT  48.83 114.69 49.16 114.54 ;
      RECT  53.09 33.82 53.44 34.17 ;
      RECT  51.25 33.33 53.85 33.62 ;
      RECT  51.76 33.82 52.11 34.17 ;
      RECT  51.45 34.48 51.74 34.64 ;
      RECT  52.59 36.99 52.88 37.28 ;
      RECT  51.25 38.45 53.85 38.74 ;
      RECT  52.17 36.45 52.46 36.74 ;
      RECT  51.43 34.33 51.76 34.48 ;
      RECT  53.09 43.38 53.44 43.03 ;
      RECT  51.25 43.87 53.85 43.58 ;
      RECT  51.76 43.38 52.11 43.03 ;
      RECT  51.45 42.72 51.74 42.56 ;
      RECT  52.59 40.21 52.88 39.92 ;
      RECT  51.25 38.75 53.85 38.46 ;
      RECT  52.17 40.75 52.46 40.46 ;
      RECT  51.43 42.87 51.76 42.72 ;
      RECT  53.09 44.08 53.44 44.43 ;
      RECT  51.25 43.59 53.85 43.88 ;
      RECT  51.76 44.08 52.11 44.43 ;
      RECT  51.45 44.74 51.74 44.9 ;
      RECT  52.59 47.25 52.88 47.54 ;
      RECT  51.25 48.71 53.85 49.0 ;
      RECT  52.17 46.71 52.46 47.0 ;
      RECT  51.43 44.59 51.76 44.74 ;
      RECT  53.09 53.64 53.44 53.29 ;
      RECT  51.25 54.13 53.85 53.84 ;
      RECT  51.76 53.64 52.11 53.29 ;
      RECT  51.45 52.98 51.74 52.82 ;
      RECT  52.59 50.47 52.88 50.18 ;
      RECT  51.25 49.01 53.85 48.72 ;
      RECT  52.17 51.01 52.46 50.72 ;
      RECT  51.43 53.13 51.76 52.98 ;
      RECT  53.09 54.34 53.44 54.69 ;
      RECT  51.25 53.85 53.85 54.14 ;
      RECT  51.76 54.34 52.11 54.69 ;
      RECT  51.45 55.0 51.74 55.16 ;
      RECT  52.59 57.51 52.88 57.8 ;
      RECT  51.25 58.97 53.85 59.26 ;
      RECT  52.17 56.97 52.46 57.26 ;
      RECT  51.43 54.85 51.76 55.0 ;
      RECT  53.09 63.9 53.44 63.55 ;
      RECT  51.25 64.39 53.85 64.1 ;
      RECT  51.76 63.9 52.11 63.55 ;
      RECT  51.45 63.24 51.74 63.08 ;
      RECT  52.59 60.73 52.88 60.44 ;
      RECT  51.25 59.27 53.85 58.98 ;
      RECT  52.17 61.27 52.46 60.98 ;
      RECT  51.43 63.39 51.76 63.24 ;
      RECT  53.09 64.6 53.44 64.95 ;
      RECT  51.25 64.11 53.85 64.4 ;
      RECT  51.76 64.6 52.11 64.95 ;
      RECT  51.45 65.26 51.74 65.42 ;
      RECT  52.59 67.77 52.88 68.06 ;
      RECT  51.25 69.23 53.85 69.52 ;
      RECT  52.17 67.23 52.46 67.52 ;
      RECT  51.43 65.11 51.76 65.26 ;
      RECT  53.09 74.16 53.44 73.81 ;
      RECT  51.25 74.65 53.85 74.36 ;
      RECT  51.76 74.16 52.11 73.81 ;
      RECT  51.45 73.5 51.74 73.34 ;
      RECT  52.59 70.99 52.88 70.7 ;
      RECT  51.25 69.53 53.85 69.24 ;
      RECT  52.17 71.53 52.46 71.24 ;
      RECT  51.43 73.65 51.76 73.5 ;
      RECT  53.09 74.86 53.44 75.21 ;
      RECT  51.25 74.37 53.85 74.66 ;
      RECT  51.76 74.86 52.11 75.21 ;
      RECT  51.45 75.52 51.74 75.68 ;
      RECT  52.59 78.03 52.88 78.32 ;
      RECT  51.25 79.49 53.85 79.78 ;
      RECT  52.17 77.49 52.46 77.78 ;
      RECT  51.43 75.37 51.76 75.52 ;
      RECT  53.09 84.42 53.44 84.07 ;
      RECT  51.25 84.91 53.85 84.62 ;
      RECT  51.76 84.42 52.11 84.07 ;
      RECT  51.45 83.76 51.74 83.6 ;
      RECT  52.59 81.25 52.88 80.96 ;
      RECT  51.25 79.79 53.85 79.5 ;
      RECT  52.17 81.79 52.46 81.5 ;
      RECT  51.43 83.91 51.76 83.76 ;
      RECT  53.09 85.12 53.44 85.47 ;
      RECT  51.25 84.63 53.85 84.92 ;
      RECT  51.76 85.12 52.11 85.47 ;
      RECT  51.45 85.78 51.74 85.94 ;
      RECT  52.59 88.29 52.88 88.58 ;
      RECT  51.25 89.75 53.85 90.04 ;
      RECT  52.17 87.75 52.46 88.04 ;
      RECT  51.43 85.63 51.76 85.78 ;
      RECT  53.09 94.68 53.44 94.33 ;
      RECT  51.25 95.17 53.85 94.88 ;
      RECT  51.76 94.68 52.11 94.33 ;
      RECT  51.45 94.02 51.74 93.86 ;
      RECT  52.59 91.51 52.88 91.22 ;
      RECT  51.25 90.05 53.85 89.76 ;
      RECT  52.17 92.05 52.46 91.76 ;
      RECT  51.43 94.17 51.76 94.02 ;
      RECT  53.09 95.38 53.44 95.73 ;
      RECT  51.25 94.89 53.85 95.18 ;
      RECT  51.76 95.38 52.11 95.73 ;
      RECT  51.45 96.04 51.74 96.2 ;
      RECT  52.59 98.55 52.88 98.84 ;
      RECT  51.25 100.01 53.85 100.3 ;
      RECT  52.17 98.01 52.46 98.3 ;
      RECT  51.43 95.89 51.76 96.04 ;
      RECT  53.09 104.94 53.44 104.59 ;
      RECT  51.25 105.43 53.85 105.14 ;
      RECT  51.76 104.94 52.11 104.59 ;
      RECT  51.45 104.28 51.74 104.12 ;
      RECT  52.59 101.77 52.88 101.48 ;
      RECT  51.25 100.31 53.85 100.02 ;
      RECT  52.17 102.31 52.46 102.02 ;
      RECT  51.43 104.43 51.76 104.28 ;
      RECT  53.09 105.64 53.44 105.99 ;
      RECT  51.25 105.15 53.85 105.44 ;
      RECT  51.76 105.64 52.11 105.99 ;
      RECT  51.45 106.3 51.74 106.46 ;
      RECT  52.59 108.81 52.88 109.1 ;
      RECT  51.25 110.27 53.85 110.56 ;
      RECT  52.17 108.27 52.46 108.56 ;
      RECT  51.43 106.15 51.76 106.3 ;
      RECT  53.09 115.2 53.44 114.85 ;
      RECT  51.25 115.69 53.85 115.4 ;
      RECT  51.76 115.2 52.11 114.85 ;
      RECT  51.45 114.54 51.74 114.38 ;
      RECT  52.59 112.03 52.88 111.74 ;
      RECT  51.25 110.57 53.85 110.28 ;
      RECT  52.17 112.57 52.46 112.28 ;
      RECT  51.43 114.69 51.76 114.54 ;
      RECT  48.65 34.48 53.85 34.64 ;
      RECT  48.65 42.56 53.85 42.72 ;
      RECT  48.65 44.74 53.85 44.9 ;
      RECT  48.65 52.82 53.85 52.98 ;
      RECT  48.65 55.0 53.85 55.16 ;
      RECT  48.65 63.08 53.85 63.24 ;
      RECT  48.65 65.26 53.85 65.42 ;
      RECT  48.65 73.34 53.85 73.5 ;
      RECT  48.65 75.52 53.85 75.68 ;
      RECT  48.65 83.6 53.85 83.76 ;
      RECT  48.65 85.78 53.85 85.94 ;
      RECT  48.65 93.86 53.85 94.02 ;
      RECT  48.65 96.04 53.85 96.2 ;
      RECT  48.65 104.12 53.85 104.28 ;
      RECT  48.65 106.3 53.85 106.46 ;
      RECT  48.65 114.38 53.85 114.54 ;
      RECT  48.65 100.01 51.25 100.3 ;
      RECT  51.25 48.72 53.85 49.01 ;
      RECT  51.25 110.28 53.85 110.57 ;
      RECT  48.65 69.24 51.25 69.53 ;
      RECT  48.65 58.97 51.25 59.26 ;
      RECT  51.25 58.97 53.85 59.26 ;
      RECT  48.65 89.75 51.25 90.04 ;
      RECT  48.65 89.76 51.25 90.05 ;
      RECT  51.25 89.75 53.85 90.04 ;
      RECT  48.65 69.23 51.25 69.52 ;
      RECT  48.65 48.71 51.25 49.0 ;
      RECT  48.65 79.49 51.25 79.78 ;
      RECT  51.25 89.76 53.85 90.05 ;
      RECT  48.65 48.72 51.25 49.01 ;
      RECT  48.65 110.27 51.25 110.56 ;
      RECT  51.25 69.24 53.85 69.53 ;
      RECT  48.65 38.46 51.25 38.75 ;
      RECT  51.25 100.02 53.85 100.31 ;
      RECT  51.25 100.01 53.85 100.3 ;
      RECT  51.25 38.46 53.85 38.75 ;
      RECT  51.25 58.98 53.85 59.27 ;
      RECT  51.25 79.5 53.85 79.79 ;
      RECT  51.25 79.49 53.85 79.78 ;
      RECT  48.65 58.98 51.25 59.27 ;
      RECT  51.25 110.27 53.85 110.56 ;
      RECT  51.25 48.71 53.85 49.0 ;
      RECT  48.65 79.5 51.25 79.79 ;
      RECT  48.65 38.45 51.25 38.74 ;
      RECT  48.65 100.02 51.25 100.31 ;
      RECT  51.25 69.23 53.85 69.52 ;
      RECT  48.65 110.28 51.25 110.57 ;
      RECT  51.25 38.45 53.85 38.74 ;
      RECT  48.65 53.84 51.25 54.13 ;
      RECT  51.25 94.88 53.85 95.17 ;
      RECT  51.25 84.62 53.85 84.91 ;
      RECT  48.65 74.36 51.25 74.65 ;
      RECT  51.25 64.1 53.85 64.39 ;
      RECT  48.65 33.33 51.25 33.62 ;
      RECT  51.25 53.85 53.85 54.14 ;
      RECT  48.65 43.59 51.25 43.88 ;
      RECT  51.25 33.33 53.85 33.62 ;
      RECT  51.25 115.4 53.85 115.69 ;
      RECT  48.65 43.58 51.25 43.87 ;
      RECT  48.65 64.11 51.25 64.4 ;
      RECT  48.65 105.15 51.25 105.44 ;
      RECT  51.25 53.84 53.85 54.13 ;
      RECT  51.25 94.89 53.85 95.18 ;
      RECT  48.65 64.1 51.25 64.39 ;
      RECT  51.25 74.37 53.85 74.66 ;
      RECT  48.65 53.85 51.25 54.14 ;
      RECT  51.25 43.58 53.85 43.87 ;
      RECT  48.65 105.14 51.25 105.43 ;
      RECT  51.25 64.11 53.85 64.4 ;
      RECT  48.65 84.63 51.25 84.92 ;
      RECT  51.25 105.14 53.85 105.43 ;
      RECT  48.65 94.88 51.25 95.17 ;
      RECT  48.65 74.37 51.25 74.66 ;
      RECT  48.65 115.4 51.25 115.69 ;
      RECT  48.65 84.62 51.25 84.91 ;
      RECT  51.25 74.36 53.85 74.65 ;
      RECT  51.25 105.15 53.85 105.44 ;
      RECT  48.65 94.89 51.25 95.18 ;
      RECT  51.25 43.59 53.85 43.88 ;
      RECT  51.25 84.63 53.85 84.92 ;
      RECT  47.89 23.56 48.24 23.91 ;
      RECT  46.05 23.07 48.65 23.36 ;
      RECT  46.56 23.56 46.91 23.91 ;
      RECT  46.25 24.22 46.54 24.38 ;
      RECT  47.39 26.73 47.68 27.02 ;
      RECT  46.05 28.19 48.65 28.48 ;
      RECT  46.97 26.19 47.26 26.48 ;
      RECT  46.23 24.07 46.56 24.22 ;
      RECT  47.89 33.12 48.24 32.77 ;
      RECT  46.05 33.61 48.65 33.32 ;
      RECT  46.56 33.12 46.91 32.77 ;
      RECT  46.25 32.46 46.54 32.3 ;
      RECT  47.39 29.95 47.68 29.66 ;
      RECT  46.05 28.49 48.65 28.2 ;
      RECT  46.97 30.49 47.26 30.2 ;
      RECT  46.23 32.61 46.56 32.46 ;
      RECT  47.89 33.82 48.24 34.17 ;
      RECT  46.05 33.33 48.65 33.62 ;
      RECT  46.56 33.82 46.91 34.17 ;
      RECT  46.25 34.48 46.54 34.64 ;
      RECT  47.39 36.99 47.68 37.28 ;
      RECT  46.05 38.45 48.65 38.74 ;
      RECT  46.97 36.45 47.26 36.74 ;
      RECT  46.23 34.33 46.56 34.48 ;
      RECT  47.89 43.38 48.24 43.03 ;
      RECT  46.05 43.87 48.65 43.58 ;
      RECT  46.56 43.38 46.91 43.03 ;
      RECT  46.25 42.72 46.54 42.56 ;
      RECT  47.39 40.21 47.68 39.92 ;
      RECT  46.05 38.75 48.65 38.46 ;
      RECT  46.97 40.75 47.26 40.46 ;
      RECT  46.23 42.87 46.56 42.72 ;
      RECT  47.89 44.08 48.24 44.43 ;
      RECT  46.05 43.59 48.65 43.88 ;
      RECT  46.56 44.08 46.91 44.43 ;
      RECT  46.25 44.74 46.54 44.9 ;
      RECT  47.39 47.25 47.68 47.54 ;
      RECT  46.05 48.71 48.65 49.0 ;
      RECT  46.97 46.71 47.26 47.0 ;
      RECT  46.23 44.59 46.56 44.74 ;
      RECT  47.89 53.64 48.24 53.29 ;
      RECT  46.05 54.13 48.65 53.84 ;
      RECT  46.56 53.64 46.91 53.29 ;
      RECT  46.25 52.98 46.54 52.82 ;
      RECT  47.39 50.47 47.68 50.18 ;
      RECT  46.05 49.01 48.65 48.72 ;
      RECT  46.97 51.01 47.26 50.72 ;
      RECT  46.23 53.13 46.56 52.98 ;
      RECT  47.89 54.34 48.24 54.69 ;
      RECT  46.05 53.85 48.65 54.14 ;
      RECT  46.56 54.34 46.91 54.69 ;
      RECT  46.25 55.0 46.54 55.16 ;
      RECT  47.39 57.51 47.68 57.8 ;
      RECT  46.05 58.97 48.65 59.26 ;
      RECT  46.97 56.97 47.26 57.26 ;
      RECT  46.23 54.85 46.56 55.0 ;
      RECT  47.89 63.9 48.24 63.55 ;
      RECT  46.05 64.39 48.65 64.1 ;
      RECT  46.56 63.9 46.91 63.55 ;
      RECT  46.25 63.24 46.54 63.08 ;
      RECT  47.39 60.73 47.68 60.44 ;
      RECT  46.05 59.27 48.65 58.98 ;
      RECT  46.97 61.27 47.26 60.98 ;
      RECT  46.23 63.39 46.56 63.24 ;
      RECT  47.89 64.6 48.24 64.95 ;
      RECT  46.05 64.11 48.65 64.4 ;
      RECT  46.56 64.6 46.91 64.95 ;
      RECT  46.25 65.26 46.54 65.42 ;
      RECT  47.39 67.77 47.68 68.06 ;
      RECT  46.05 69.23 48.65 69.52 ;
      RECT  46.97 67.23 47.26 67.52 ;
      RECT  46.23 65.11 46.56 65.26 ;
      RECT  47.89 74.16 48.24 73.81 ;
      RECT  46.05 74.65 48.65 74.36 ;
      RECT  46.56 74.16 46.91 73.81 ;
      RECT  46.25 73.5 46.54 73.34 ;
      RECT  47.39 70.99 47.68 70.7 ;
      RECT  46.05 69.53 48.65 69.24 ;
      RECT  46.97 71.53 47.26 71.24 ;
      RECT  46.23 73.65 46.56 73.5 ;
      RECT  47.89 74.86 48.24 75.21 ;
      RECT  46.05 74.37 48.65 74.66 ;
      RECT  46.56 74.86 46.91 75.21 ;
      RECT  46.25 75.52 46.54 75.68 ;
      RECT  47.39 78.03 47.68 78.32 ;
      RECT  46.05 79.49 48.65 79.78 ;
      RECT  46.97 77.49 47.26 77.78 ;
      RECT  46.23 75.37 46.56 75.52 ;
      RECT  47.89 84.42 48.24 84.07 ;
      RECT  46.05 84.91 48.65 84.62 ;
      RECT  46.56 84.42 46.91 84.07 ;
      RECT  46.25 83.76 46.54 83.6 ;
      RECT  47.39 81.25 47.68 80.96 ;
      RECT  46.05 79.79 48.65 79.5 ;
      RECT  46.97 81.79 47.26 81.5 ;
      RECT  46.23 83.91 46.56 83.76 ;
      RECT  47.89 85.12 48.24 85.47 ;
      RECT  46.05 84.63 48.65 84.92 ;
      RECT  46.56 85.12 46.91 85.47 ;
      RECT  46.25 85.78 46.54 85.94 ;
      RECT  47.39 88.29 47.68 88.58 ;
      RECT  46.05 89.75 48.65 90.04 ;
      RECT  46.97 87.75 47.26 88.04 ;
      RECT  46.23 85.63 46.56 85.78 ;
      RECT  47.89 94.68 48.24 94.33 ;
      RECT  46.05 95.17 48.65 94.88 ;
      RECT  46.56 94.68 46.91 94.33 ;
      RECT  46.25 94.02 46.54 93.86 ;
      RECT  47.39 91.51 47.68 91.22 ;
      RECT  46.05 90.05 48.65 89.76 ;
      RECT  46.97 92.05 47.26 91.76 ;
      RECT  46.23 94.17 46.56 94.02 ;
      RECT  47.89 95.38 48.24 95.73 ;
      RECT  46.05 94.89 48.65 95.18 ;
      RECT  46.56 95.38 46.91 95.73 ;
      RECT  46.25 96.04 46.54 96.2 ;
      RECT  47.39 98.55 47.68 98.84 ;
      RECT  46.05 100.01 48.65 100.3 ;
      RECT  46.97 98.01 47.26 98.3 ;
      RECT  46.23 95.89 46.56 96.04 ;
      RECT  47.89 104.94 48.24 104.59 ;
      RECT  46.05 105.43 48.65 105.14 ;
      RECT  46.56 104.94 46.91 104.59 ;
      RECT  46.25 104.28 46.54 104.12 ;
      RECT  47.39 101.77 47.68 101.48 ;
      RECT  46.05 100.31 48.65 100.02 ;
      RECT  46.97 102.31 47.26 102.02 ;
      RECT  46.23 104.43 46.56 104.28 ;
      RECT  47.89 105.64 48.24 105.99 ;
      RECT  46.05 105.15 48.65 105.44 ;
      RECT  46.56 105.64 46.91 105.99 ;
      RECT  46.25 106.3 46.54 106.46 ;
      RECT  47.39 108.81 47.68 109.1 ;
      RECT  46.05 110.27 48.65 110.56 ;
      RECT  46.97 108.27 47.26 108.56 ;
      RECT  46.23 106.15 46.56 106.3 ;
      RECT  47.89 115.2 48.24 114.85 ;
      RECT  46.05 115.69 48.65 115.4 ;
      RECT  46.56 115.2 46.91 114.85 ;
      RECT  46.25 114.54 46.54 114.38 ;
      RECT  47.39 112.03 47.68 111.74 ;
      RECT  46.05 110.57 48.65 110.28 ;
      RECT  46.97 112.57 47.26 112.28 ;
      RECT  46.23 114.69 46.56 114.54 ;
      RECT  47.89 115.9 48.24 116.25 ;
      RECT  46.05 115.41 48.65 115.7 ;
      RECT  46.56 115.9 46.91 116.25 ;
      RECT  46.25 116.56 46.54 116.72 ;
      RECT  47.39 119.07 47.68 119.36 ;
      RECT  46.05 120.53 48.65 120.82 ;
      RECT  46.97 118.53 47.26 118.82 ;
      RECT  46.23 116.41 46.56 116.56 ;
      RECT  46.05 24.22 48.65 24.38 ;
      RECT  46.05 32.3 48.65 32.46 ;
      RECT  46.05 34.48 48.65 34.64 ;
      RECT  46.05 42.56 48.65 42.72 ;
      RECT  46.05 44.74 48.65 44.9 ;
      RECT  46.05 52.82 48.65 52.98 ;
      RECT  46.05 55.0 48.65 55.16 ;
      RECT  46.05 63.08 48.65 63.24 ;
      RECT  46.05 65.26 48.65 65.42 ;
      RECT  46.05 73.34 48.65 73.5 ;
      RECT  46.05 75.52 48.65 75.68 ;
      RECT  46.05 83.6 48.65 83.76 ;
      RECT  46.05 85.78 48.65 85.94 ;
      RECT  46.05 93.86 48.65 94.02 ;
      RECT  46.05 96.04 48.65 96.2 ;
      RECT  46.05 104.12 48.65 104.28 ;
      RECT  46.05 106.3 48.65 106.46 ;
      RECT  46.05 114.38 48.65 114.54 ;
      RECT  46.05 116.56 48.65 116.72 ;
      RECT  46.05 89.75 48.65 90.04 ;
      RECT  46.05 58.98 48.65 59.27 ;
      RECT  46.05 48.71 48.65 49.0 ;
      RECT  46.05 79.49 48.65 79.78 ;
      RECT  46.05 79.5 48.65 79.79 ;
      RECT  46.05 58.97 48.65 59.26 ;
      RECT  46.05 38.45 48.65 38.74 ;
      RECT  46.05 69.23 48.65 69.52 ;
      RECT  46.05 110.27 48.65 110.56 ;
      RECT  46.05 110.28 48.65 110.57 ;
      RECT  46.05 38.46 48.65 38.75 ;
      RECT  46.05 100.01 48.65 100.3 ;
      RECT  46.05 28.2 48.65 28.49 ;
      RECT  46.05 48.72 48.65 49.01 ;
      RECT  46.05 69.24 48.65 69.53 ;
      RECT  46.05 89.76 48.65 90.05 ;
      RECT  46.05 100.02 48.65 100.31 ;
      RECT  46.05 43.58 48.65 43.87 ;
      RECT  46.05 64.1 48.65 64.39 ;
      RECT  46.05 115.4 48.65 115.69 ;
      RECT  46.05 33.33 48.65 33.62 ;
      RECT  46.05 33.32 48.65 33.61 ;
      RECT  46.05 53.85 48.65 54.14 ;
      RECT  46.05 94.89 48.65 95.18 ;
      RECT  46.05 53.84 48.65 54.13 ;
      RECT  46.05 43.59 48.65 43.88 ;
      RECT  46.05 105.15 48.65 105.44 ;
      RECT  46.05 94.88 48.65 95.17 ;
      RECT  46.05 74.37 48.65 74.66 ;
      RECT  46.05 84.62 48.65 84.91 ;
      RECT  46.05 64.11 48.65 64.4 ;
      RECT  46.05 105.14 48.65 105.43 ;
      RECT  46.05 74.36 48.65 74.65 ;
      RECT  46.05 84.63 48.65 84.92 ;
      RECT  50.49 33.12 50.84 32.77 ;
      RECT  48.65 33.61 51.25 33.32 ;
      RECT  49.16 33.12 49.51 32.77 ;
      RECT  48.85 32.46 49.14 32.3 ;
      RECT  49.99 29.95 50.28 29.66 ;
      RECT  48.65 28.49 51.25 28.2 ;
      RECT  49.57 30.49 49.86 30.2 ;
      RECT  48.83 32.61 49.16 32.46 ;
      RECT  53.09 33.12 53.44 32.77 ;
      RECT  51.25 33.61 53.85 33.32 ;
      RECT  51.76 33.12 52.11 32.77 ;
      RECT  51.45 32.46 51.74 32.3 ;
      RECT  52.59 29.95 52.88 29.66 ;
      RECT  51.25 28.49 53.85 28.2 ;
      RECT  52.17 30.49 52.46 30.2 ;
      RECT  51.43 32.61 51.76 32.46 ;
      RECT  48.65 32.46 53.85 32.3 ;
      RECT  48.65 28.49 51.25 28.2 ;
      RECT  51.25 28.49 53.85 28.2 ;
      RECT  48.65 33.61 51.25 33.32 ;
      RECT  51.25 33.61 53.85 33.32 ;
      RECT  50.49 23.56 50.84 23.91 ;
      RECT  48.65 23.07 51.25 23.36 ;
      RECT  49.16 23.56 49.51 23.91 ;
      RECT  48.85 24.22 49.14 24.38 ;
      RECT  49.99 26.73 50.28 27.02 ;
      RECT  48.65 28.19 51.25 28.48 ;
      RECT  49.57 26.19 49.86 26.48 ;
      RECT  48.83 24.07 49.16 24.22 ;
      RECT  53.09 23.56 53.44 23.91 ;
      RECT  51.25 23.07 53.85 23.36 ;
      RECT  51.76 23.56 52.11 23.91 ;
      RECT  51.45 24.22 51.74 24.38 ;
      RECT  52.59 26.73 52.88 27.02 ;
      RECT  51.25 28.19 53.85 28.48 ;
      RECT  52.17 26.19 52.46 26.48 ;
      RECT  51.43 24.07 51.76 24.22 ;
      RECT  48.65 24.22 53.85 24.38 ;
      RECT  48.65 28.19 51.25 28.48 ;
      RECT  51.25 28.19 53.85 28.48 ;
      RECT  48.65 23.07 51.25 23.36 ;
      RECT  51.25 23.07 53.85 23.36 ;
      RECT  50.49 115.9 50.84 116.25 ;
      RECT  48.65 115.41 51.25 115.7 ;
      RECT  49.16 115.9 49.51 116.25 ;
      RECT  48.85 116.56 49.14 116.72 ;
      RECT  49.99 119.07 50.28 119.36 ;
      RECT  48.65 120.53 51.25 120.82 ;
      RECT  49.57 118.53 49.86 118.82 ;
      RECT  48.83 116.41 49.16 116.56 ;
      RECT  53.09 115.9 53.44 116.25 ;
      RECT  51.25 115.41 53.85 115.7 ;
      RECT  51.76 115.9 52.11 116.25 ;
      RECT  51.45 116.56 51.74 116.72 ;
      RECT  52.59 119.07 52.88 119.36 ;
      RECT  51.25 120.53 53.85 120.82 ;
      RECT  52.17 118.53 52.46 118.82 ;
      RECT  51.43 116.41 51.76 116.56 ;
      RECT  48.65 116.56 53.85 116.72 ;
      RECT  48.65 120.53 51.25 120.82 ;
      RECT  51.25 120.53 53.85 120.82 ;
      RECT  48.65 115.41 51.25 115.7 ;
      RECT  51.25 115.41 53.85 115.7 ;
      RECT  45.29 23.56 45.64 23.91 ;
      RECT  43.45 23.07 46.05 23.36 ;
      RECT  43.96 23.56 44.31 23.91 ;
      RECT  43.65 24.22 43.94 24.38 ;
      RECT  44.79 26.73 45.08 27.02 ;
      RECT  43.45 28.19 46.05 28.48 ;
      RECT  44.37 26.19 44.66 26.48 ;
      RECT  43.63 24.07 43.96 24.22 ;
      RECT  45.29 33.12 45.64 32.77 ;
      RECT  43.45 33.61 46.05 33.32 ;
      RECT  43.96 33.12 44.31 32.77 ;
      RECT  43.65 32.46 43.94 32.3 ;
      RECT  44.79 29.95 45.08 29.66 ;
      RECT  43.45 28.49 46.05 28.2 ;
      RECT  44.37 30.49 44.66 30.2 ;
      RECT  43.63 32.61 43.96 32.46 ;
      RECT  45.29 33.82 45.64 34.17 ;
      RECT  43.45 33.33 46.05 33.62 ;
      RECT  43.96 33.82 44.31 34.17 ;
      RECT  43.65 34.48 43.94 34.64 ;
      RECT  44.79 36.99 45.08 37.28 ;
      RECT  43.45 38.45 46.05 38.74 ;
      RECT  44.37 36.45 44.66 36.74 ;
      RECT  43.63 34.33 43.96 34.48 ;
      RECT  45.29 43.38 45.64 43.03 ;
      RECT  43.45 43.87 46.05 43.58 ;
      RECT  43.96 43.38 44.31 43.03 ;
      RECT  43.65 42.72 43.94 42.56 ;
      RECT  44.79 40.21 45.08 39.92 ;
      RECT  43.45 38.75 46.05 38.46 ;
      RECT  44.37 40.75 44.66 40.46 ;
      RECT  43.63 42.87 43.96 42.72 ;
      RECT  45.29 44.08 45.64 44.43 ;
      RECT  43.45 43.59 46.05 43.88 ;
      RECT  43.96 44.08 44.31 44.43 ;
      RECT  43.65 44.74 43.94 44.9 ;
      RECT  44.79 47.25 45.08 47.54 ;
      RECT  43.45 48.71 46.05 49.0 ;
      RECT  44.37 46.71 44.66 47.0 ;
      RECT  43.63 44.59 43.96 44.74 ;
      RECT  45.29 53.64 45.64 53.29 ;
      RECT  43.45 54.13 46.05 53.84 ;
      RECT  43.96 53.64 44.31 53.29 ;
      RECT  43.65 52.98 43.94 52.82 ;
      RECT  44.79 50.47 45.08 50.18 ;
      RECT  43.45 49.01 46.05 48.72 ;
      RECT  44.37 51.01 44.66 50.72 ;
      RECT  43.63 53.13 43.96 52.98 ;
      RECT  45.29 54.34 45.64 54.69 ;
      RECT  43.45 53.85 46.05 54.14 ;
      RECT  43.96 54.34 44.31 54.69 ;
      RECT  43.65 55.0 43.94 55.16 ;
      RECT  44.79 57.51 45.08 57.8 ;
      RECT  43.45 58.97 46.05 59.26 ;
      RECT  44.37 56.97 44.66 57.26 ;
      RECT  43.63 54.85 43.96 55.0 ;
      RECT  45.29 63.9 45.64 63.55 ;
      RECT  43.45 64.39 46.05 64.1 ;
      RECT  43.96 63.9 44.31 63.55 ;
      RECT  43.65 63.24 43.94 63.08 ;
      RECT  44.79 60.73 45.08 60.44 ;
      RECT  43.45 59.27 46.05 58.98 ;
      RECT  44.37 61.27 44.66 60.98 ;
      RECT  43.63 63.39 43.96 63.24 ;
      RECT  45.29 64.6 45.64 64.95 ;
      RECT  43.45 64.11 46.05 64.4 ;
      RECT  43.96 64.6 44.31 64.95 ;
      RECT  43.65 65.26 43.94 65.42 ;
      RECT  44.79 67.77 45.08 68.06 ;
      RECT  43.45 69.23 46.05 69.52 ;
      RECT  44.37 67.23 44.66 67.52 ;
      RECT  43.63 65.11 43.96 65.26 ;
      RECT  45.29 74.16 45.64 73.81 ;
      RECT  43.45 74.65 46.05 74.36 ;
      RECT  43.96 74.16 44.31 73.81 ;
      RECT  43.65 73.5 43.94 73.34 ;
      RECT  44.79 70.99 45.08 70.7 ;
      RECT  43.45 69.53 46.05 69.24 ;
      RECT  44.37 71.53 44.66 71.24 ;
      RECT  43.63 73.65 43.96 73.5 ;
      RECT  45.29 74.86 45.64 75.21 ;
      RECT  43.45 74.37 46.05 74.66 ;
      RECT  43.96 74.86 44.31 75.21 ;
      RECT  43.65 75.52 43.94 75.68 ;
      RECT  44.79 78.03 45.08 78.32 ;
      RECT  43.45 79.49 46.05 79.78 ;
      RECT  44.37 77.49 44.66 77.78 ;
      RECT  43.63 75.37 43.96 75.52 ;
      RECT  45.29 84.42 45.64 84.07 ;
      RECT  43.45 84.91 46.05 84.62 ;
      RECT  43.96 84.42 44.31 84.07 ;
      RECT  43.65 83.76 43.94 83.6 ;
      RECT  44.79 81.25 45.08 80.96 ;
      RECT  43.45 79.79 46.05 79.5 ;
      RECT  44.37 81.79 44.66 81.5 ;
      RECT  43.63 83.91 43.96 83.76 ;
      RECT  45.29 85.12 45.64 85.47 ;
      RECT  43.45 84.63 46.05 84.92 ;
      RECT  43.96 85.12 44.31 85.47 ;
      RECT  43.65 85.78 43.94 85.94 ;
      RECT  44.79 88.29 45.08 88.58 ;
      RECT  43.45 89.75 46.05 90.04 ;
      RECT  44.37 87.75 44.66 88.04 ;
      RECT  43.63 85.63 43.96 85.78 ;
      RECT  45.29 94.68 45.64 94.33 ;
      RECT  43.45 95.17 46.05 94.88 ;
      RECT  43.96 94.68 44.31 94.33 ;
      RECT  43.65 94.02 43.94 93.86 ;
      RECT  44.79 91.51 45.08 91.22 ;
      RECT  43.45 90.05 46.05 89.76 ;
      RECT  44.37 92.05 44.66 91.76 ;
      RECT  43.63 94.17 43.96 94.02 ;
      RECT  45.29 95.38 45.64 95.73 ;
      RECT  43.45 94.89 46.05 95.18 ;
      RECT  43.96 95.38 44.31 95.73 ;
      RECT  43.65 96.04 43.94 96.2 ;
      RECT  44.79 98.55 45.08 98.84 ;
      RECT  43.45 100.01 46.05 100.3 ;
      RECT  44.37 98.01 44.66 98.3 ;
      RECT  43.63 95.89 43.96 96.04 ;
      RECT  45.29 104.94 45.64 104.59 ;
      RECT  43.45 105.43 46.05 105.14 ;
      RECT  43.96 104.94 44.31 104.59 ;
      RECT  43.65 104.28 43.94 104.12 ;
      RECT  44.79 101.77 45.08 101.48 ;
      RECT  43.45 100.31 46.05 100.02 ;
      RECT  44.37 102.31 44.66 102.02 ;
      RECT  43.63 104.43 43.96 104.28 ;
      RECT  45.29 105.64 45.64 105.99 ;
      RECT  43.45 105.15 46.05 105.44 ;
      RECT  43.96 105.64 44.31 105.99 ;
      RECT  43.65 106.3 43.94 106.46 ;
      RECT  44.79 108.81 45.08 109.1 ;
      RECT  43.45 110.27 46.05 110.56 ;
      RECT  44.37 108.27 44.66 108.56 ;
      RECT  43.63 106.15 43.96 106.3 ;
      RECT  45.29 115.2 45.64 114.85 ;
      RECT  43.45 115.69 46.05 115.4 ;
      RECT  43.96 115.2 44.31 114.85 ;
      RECT  43.65 114.54 43.94 114.38 ;
      RECT  44.79 112.03 45.08 111.74 ;
      RECT  43.45 110.57 46.05 110.28 ;
      RECT  44.37 112.57 44.66 112.28 ;
      RECT  43.63 114.69 43.96 114.54 ;
      RECT  45.29 115.9 45.64 116.25 ;
      RECT  43.45 115.41 46.05 115.7 ;
      RECT  43.96 115.9 44.31 116.25 ;
      RECT  43.65 116.56 43.94 116.72 ;
      RECT  44.79 119.07 45.08 119.36 ;
      RECT  43.45 120.53 46.05 120.82 ;
      RECT  44.37 118.53 44.66 118.82 ;
      RECT  43.63 116.41 43.96 116.56 ;
      RECT  43.45 24.22 46.05 24.38 ;
      RECT  43.45 32.3 46.05 32.46 ;
      RECT  43.45 34.48 46.05 34.64 ;
      RECT  43.45 42.56 46.05 42.72 ;
      RECT  43.45 44.74 46.05 44.9 ;
      RECT  43.45 52.82 46.05 52.98 ;
      RECT  43.45 55.0 46.05 55.16 ;
      RECT  43.45 63.08 46.05 63.24 ;
      RECT  43.45 65.26 46.05 65.42 ;
      RECT  43.45 73.34 46.05 73.5 ;
      RECT  43.45 75.52 46.05 75.68 ;
      RECT  43.45 83.6 46.05 83.76 ;
      RECT  43.45 85.78 46.05 85.94 ;
      RECT  43.45 93.86 46.05 94.02 ;
      RECT  43.45 96.04 46.05 96.2 ;
      RECT  43.45 104.12 46.05 104.28 ;
      RECT  43.45 106.3 46.05 106.46 ;
      RECT  43.45 114.38 46.05 114.54 ;
      RECT  43.45 116.56 46.05 116.72 ;
      RECT  43.45 89.75 46.05 90.04 ;
      RECT  43.45 58.98 46.05 59.27 ;
      RECT  43.45 48.71 46.05 49.0 ;
      RECT  43.45 79.49 46.05 79.78 ;
      RECT  43.45 79.5 46.05 79.79 ;
      RECT  43.45 58.97 46.05 59.26 ;
      RECT  43.45 38.45 46.05 38.74 ;
      RECT  43.45 69.23 46.05 69.52 ;
      RECT  43.45 110.27 46.05 110.56 ;
      RECT  43.45 110.28 46.05 110.57 ;
      RECT  43.45 38.46 46.05 38.75 ;
      RECT  43.45 100.01 46.05 100.3 ;
      RECT  43.45 28.2 46.05 28.49 ;
      RECT  43.45 48.72 46.05 49.01 ;
      RECT  43.45 120.53 46.05 120.82 ;
      RECT  43.45 69.24 46.05 69.53 ;
      RECT  43.45 28.19 46.05 28.48 ;
      RECT  43.45 89.76 46.05 90.05 ;
      RECT  43.45 100.02 46.05 100.31 ;
      RECT  43.45 43.58 46.05 43.87 ;
      RECT  43.45 64.1 46.05 64.39 ;
      RECT  43.45 23.07 46.05 23.36 ;
      RECT  43.45 115.4 46.05 115.69 ;
      RECT  43.45 33.33 46.05 33.62 ;
      RECT  43.45 33.32 46.05 33.61 ;
      RECT  43.45 53.85 46.05 54.14 ;
      RECT  43.45 94.89 46.05 95.18 ;
      RECT  43.45 115.41 46.05 115.7 ;
      RECT  43.45 53.84 46.05 54.13 ;
      RECT  43.45 43.59 46.05 43.88 ;
      RECT  43.45 105.15 46.05 105.44 ;
      RECT  43.45 94.88 46.05 95.17 ;
      RECT  43.45 74.37 46.05 74.66 ;
      RECT  43.45 84.62 46.05 84.91 ;
      RECT  43.45 64.11 46.05 64.4 ;
      RECT  43.45 105.14 46.05 105.43 ;
      RECT  43.45 74.36 46.05 74.65 ;
      RECT  43.45 84.63 46.05 84.92 ;
      RECT  55.69 23.56 56.04 23.91 ;
      RECT  53.85 23.07 56.45 23.36 ;
      RECT  54.36 23.56 54.71 23.91 ;
      RECT  54.05 24.22 54.34 24.38 ;
      RECT  55.19 26.73 55.48 27.02 ;
      RECT  53.85 28.19 56.45 28.48 ;
      RECT  54.77 26.19 55.06 26.48 ;
      RECT  54.03 24.07 54.36 24.22 ;
      RECT  55.69 33.12 56.04 32.77 ;
      RECT  53.85 33.61 56.45 33.32 ;
      RECT  54.36 33.12 54.71 32.77 ;
      RECT  54.05 32.46 54.34 32.3 ;
      RECT  55.19 29.95 55.48 29.66 ;
      RECT  53.85 28.49 56.45 28.2 ;
      RECT  54.77 30.49 55.06 30.2 ;
      RECT  54.03 32.61 54.36 32.46 ;
      RECT  55.69 33.82 56.04 34.17 ;
      RECT  53.85 33.33 56.45 33.62 ;
      RECT  54.36 33.82 54.71 34.17 ;
      RECT  54.05 34.48 54.34 34.64 ;
      RECT  55.19 36.99 55.48 37.28 ;
      RECT  53.85 38.45 56.45 38.74 ;
      RECT  54.77 36.45 55.06 36.74 ;
      RECT  54.03 34.33 54.36 34.48 ;
      RECT  55.69 43.38 56.04 43.03 ;
      RECT  53.85 43.87 56.45 43.58 ;
      RECT  54.36 43.38 54.71 43.03 ;
      RECT  54.05 42.72 54.34 42.56 ;
      RECT  55.19 40.21 55.48 39.92 ;
      RECT  53.85 38.75 56.45 38.46 ;
      RECT  54.77 40.75 55.06 40.46 ;
      RECT  54.03 42.87 54.36 42.72 ;
      RECT  55.69 44.08 56.04 44.43 ;
      RECT  53.85 43.59 56.45 43.88 ;
      RECT  54.36 44.08 54.71 44.43 ;
      RECT  54.05 44.74 54.34 44.9 ;
      RECT  55.19 47.25 55.48 47.54 ;
      RECT  53.85 48.71 56.45 49.0 ;
      RECT  54.77 46.71 55.06 47.0 ;
      RECT  54.03 44.59 54.36 44.74 ;
      RECT  55.69 53.64 56.04 53.29 ;
      RECT  53.85 54.13 56.45 53.84 ;
      RECT  54.36 53.64 54.71 53.29 ;
      RECT  54.05 52.98 54.34 52.82 ;
      RECT  55.19 50.47 55.48 50.18 ;
      RECT  53.85 49.01 56.45 48.72 ;
      RECT  54.77 51.01 55.06 50.72 ;
      RECT  54.03 53.13 54.36 52.98 ;
      RECT  55.69 54.34 56.04 54.69 ;
      RECT  53.85 53.85 56.45 54.14 ;
      RECT  54.36 54.34 54.71 54.69 ;
      RECT  54.05 55.0 54.34 55.16 ;
      RECT  55.19 57.51 55.48 57.8 ;
      RECT  53.85 58.97 56.45 59.26 ;
      RECT  54.77 56.97 55.06 57.26 ;
      RECT  54.03 54.85 54.36 55.0 ;
      RECT  55.69 63.9 56.04 63.55 ;
      RECT  53.85 64.39 56.45 64.1 ;
      RECT  54.36 63.9 54.71 63.55 ;
      RECT  54.05 63.24 54.34 63.08 ;
      RECT  55.19 60.73 55.48 60.44 ;
      RECT  53.85 59.27 56.45 58.98 ;
      RECT  54.77 61.27 55.06 60.98 ;
      RECT  54.03 63.39 54.36 63.24 ;
      RECT  55.69 64.6 56.04 64.95 ;
      RECT  53.85 64.11 56.45 64.4 ;
      RECT  54.36 64.6 54.71 64.95 ;
      RECT  54.05 65.26 54.34 65.42 ;
      RECT  55.19 67.77 55.48 68.06 ;
      RECT  53.85 69.23 56.45 69.52 ;
      RECT  54.77 67.23 55.06 67.52 ;
      RECT  54.03 65.11 54.36 65.26 ;
      RECT  55.69 74.16 56.04 73.81 ;
      RECT  53.85 74.65 56.45 74.36 ;
      RECT  54.36 74.16 54.71 73.81 ;
      RECT  54.05 73.5 54.34 73.34 ;
      RECT  55.19 70.99 55.48 70.7 ;
      RECT  53.85 69.53 56.45 69.24 ;
      RECT  54.77 71.53 55.06 71.24 ;
      RECT  54.03 73.65 54.36 73.5 ;
      RECT  55.69 74.86 56.04 75.21 ;
      RECT  53.85 74.37 56.45 74.66 ;
      RECT  54.36 74.86 54.71 75.21 ;
      RECT  54.05 75.52 54.34 75.68 ;
      RECT  55.19 78.03 55.48 78.32 ;
      RECT  53.85 79.49 56.45 79.78 ;
      RECT  54.77 77.49 55.06 77.78 ;
      RECT  54.03 75.37 54.36 75.52 ;
      RECT  55.69 84.42 56.04 84.07 ;
      RECT  53.85 84.91 56.45 84.62 ;
      RECT  54.36 84.42 54.71 84.07 ;
      RECT  54.05 83.76 54.34 83.6 ;
      RECT  55.19 81.25 55.48 80.96 ;
      RECT  53.85 79.79 56.45 79.5 ;
      RECT  54.77 81.79 55.06 81.5 ;
      RECT  54.03 83.91 54.36 83.76 ;
      RECT  55.69 85.12 56.04 85.47 ;
      RECT  53.85 84.63 56.45 84.92 ;
      RECT  54.36 85.12 54.71 85.47 ;
      RECT  54.05 85.78 54.34 85.94 ;
      RECT  55.19 88.29 55.48 88.58 ;
      RECT  53.85 89.75 56.45 90.04 ;
      RECT  54.77 87.75 55.06 88.04 ;
      RECT  54.03 85.63 54.36 85.78 ;
      RECT  55.69 94.68 56.04 94.33 ;
      RECT  53.85 95.17 56.45 94.88 ;
      RECT  54.36 94.68 54.71 94.33 ;
      RECT  54.05 94.02 54.34 93.86 ;
      RECT  55.19 91.51 55.48 91.22 ;
      RECT  53.85 90.05 56.45 89.76 ;
      RECT  54.77 92.05 55.06 91.76 ;
      RECT  54.03 94.17 54.36 94.02 ;
      RECT  55.69 95.38 56.04 95.73 ;
      RECT  53.85 94.89 56.45 95.18 ;
      RECT  54.36 95.38 54.71 95.73 ;
      RECT  54.05 96.04 54.34 96.2 ;
      RECT  55.19 98.55 55.48 98.84 ;
      RECT  53.85 100.01 56.45 100.3 ;
      RECT  54.77 98.01 55.06 98.3 ;
      RECT  54.03 95.89 54.36 96.04 ;
      RECT  55.69 104.94 56.04 104.59 ;
      RECT  53.85 105.43 56.45 105.14 ;
      RECT  54.36 104.94 54.71 104.59 ;
      RECT  54.05 104.28 54.34 104.12 ;
      RECT  55.19 101.77 55.48 101.48 ;
      RECT  53.85 100.31 56.45 100.02 ;
      RECT  54.77 102.31 55.06 102.02 ;
      RECT  54.03 104.43 54.36 104.28 ;
      RECT  55.69 105.64 56.04 105.99 ;
      RECT  53.85 105.15 56.45 105.44 ;
      RECT  54.36 105.64 54.71 105.99 ;
      RECT  54.05 106.3 54.34 106.46 ;
      RECT  55.19 108.81 55.48 109.1 ;
      RECT  53.85 110.27 56.45 110.56 ;
      RECT  54.77 108.27 55.06 108.56 ;
      RECT  54.03 106.15 54.36 106.3 ;
      RECT  55.69 115.2 56.04 114.85 ;
      RECT  53.85 115.69 56.45 115.4 ;
      RECT  54.36 115.2 54.71 114.85 ;
      RECT  54.05 114.54 54.34 114.38 ;
      RECT  55.19 112.03 55.48 111.74 ;
      RECT  53.85 110.57 56.45 110.28 ;
      RECT  54.77 112.57 55.06 112.28 ;
      RECT  54.03 114.69 54.36 114.54 ;
      RECT  55.69 115.9 56.04 116.25 ;
      RECT  53.85 115.41 56.45 115.7 ;
      RECT  54.36 115.9 54.71 116.25 ;
      RECT  54.05 116.56 54.34 116.72 ;
      RECT  55.19 119.07 55.48 119.36 ;
      RECT  53.85 120.53 56.45 120.82 ;
      RECT  54.77 118.53 55.06 118.82 ;
      RECT  54.03 116.41 54.36 116.56 ;
      RECT  53.85 24.22 56.45 24.38 ;
      RECT  53.85 32.3 56.45 32.46 ;
      RECT  53.85 34.48 56.45 34.64 ;
      RECT  53.85 42.56 56.45 42.72 ;
      RECT  53.85 44.74 56.45 44.9 ;
      RECT  53.85 52.82 56.45 52.98 ;
      RECT  53.85 55.0 56.45 55.16 ;
      RECT  53.85 63.08 56.45 63.24 ;
      RECT  53.85 65.26 56.45 65.42 ;
      RECT  53.85 73.34 56.45 73.5 ;
      RECT  53.85 75.52 56.45 75.68 ;
      RECT  53.85 83.6 56.45 83.76 ;
      RECT  53.85 85.78 56.45 85.94 ;
      RECT  53.85 93.86 56.45 94.02 ;
      RECT  53.85 96.04 56.45 96.2 ;
      RECT  53.85 104.12 56.45 104.28 ;
      RECT  53.85 106.3 56.45 106.46 ;
      RECT  53.85 114.38 56.45 114.54 ;
      RECT  53.85 116.56 56.45 116.72 ;
      RECT  53.85 89.75 56.45 90.04 ;
      RECT  53.85 58.98 56.45 59.27 ;
      RECT  53.85 48.71 56.45 49.0 ;
      RECT  53.85 79.49 56.45 79.78 ;
      RECT  53.85 79.5 56.45 79.79 ;
      RECT  53.85 58.97 56.45 59.26 ;
      RECT  53.85 38.45 56.45 38.74 ;
      RECT  53.85 69.23 56.45 69.52 ;
      RECT  53.85 110.27 56.45 110.56 ;
      RECT  53.85 110.28 56.45 110.57 ;
      RECT  53.85 38.46 56.45 38.75 ;
      RECT  53.85 100.01 56.45 100.3 ;
      RECT  53.85 28.2 56.45 28.49 ;
      RECT  53.85 48.72 56.45 49.01 ;
      RECT  53.85 120.53 56.45 120.82 ;
      RECT  53.85 69.24 56.45 69.53 ;
      RECT  53.85 28.19 56.45 28.48 ;
      RECT  53.85 89.76 56.45 90.05 ;
      RECT  53.85 100.02 56.45 100.31 ;
      RECT  53.85 43.58 56.45 43.87 ;
      RECT  53.85 64.1 56.45 64.39 ;
      RECT  53.85 23.07 56.45 23.36 ;
      RECT  53.85 115.4 56.45 115.69 ;
      RECT  53.85 33.33 56.45 33.62 ;
      RECT  53.85 33.32 56.45 33.61 ;
      RECT  53.85 53.85 56.45 54.14 ;
      RECT  53.85 94.89 56.45 95.18 ;
      RECT  53.85 115.41 56.45 115.7 ;
      RECT  53.85 53.84 56.45 54.13 ;
      RECT  53.85 43.59 56.45 43.88 ;
      RECT  53.85 105.15 56.45 105.44 ;
      RECT  53.85 94.88 56.45 95.17 ;
      RECT  53.85 74.37 56.45 74.66 ;
      RECT  53.85 84.62 56.45 84.91 ;
      RECT  53.85 64.11 56.45 64.4 ;
      RECT  53.85 105.14 56.45 105.43 ;
      RECT  53.85 74.36 56.45 74.65 ;
      RECT  53.85 84.63 56.45 84.92 ;
      RECT  42.55 32.3 57.35 32.46 ;
      RECT  42.55 34.48 57.35 34.64 ;
      RECT  42.55 42.56 57.35 42.72 ;
      RECT  42.55 44.74 57.35 44.9 ;
      RECT  42.55 52.82 57.35 52.98 ;
      RECT  42.55 55.0 57.35 55.16 ;
      RECT  42.55 63.08 57.35 63.24 ;
      RECT  42.55 65.26 57.35 65.42 ;
      RECT  42.55 73.34 57.35 73.5 ;
      RECT  42.55 75.52 57.35 75.68 ;
      RECT  42.55 83.6 57.35 83.76 ;
      RECT  42.55 85.78 57.35 85.94 ;
      RECT  42.55 93.86 57.35 94.02 ;
      RECT  42.55 96.04 57.35 96.2 ;
      RECT  42.55 104.12 57.35 104.28 ;
      RECT  42.55 106.3 57.35 106.46 ;
      RECT  42.55 114.38 57.35 114.54 ;
      RECT  46.05 79.5 48.65 79.79 ;
      RECT  46.05 58.97 48.65 59.26 ;
      RECT  46.05 48.71 48.65 49.0 ;
      RECT  46.05 110.28 48.65 110.57 ;
      RECT  46.05 38.46 48.65 38.75 ;
      RECT  46.05 110.27 48.65 110.56 ;
      RECT  46.05 69.24 48.65 69.53 ;
      RECT  46.05 69.23 48.65 69.52 ;
      RECT  46.05 100.01 48.65 100.3 ;
      RECT  46.05 58.98 48.65 59.27 ;
      RECT  46.05 89.76 48.65 90.05 ;
      RECT  46.05 79.49 48.65 79.78 ;
      RECT  46.05 38.45 48.65 38.74 ;
      RECT  46.05 48.72 48.65 49.01 ;
      RECT  46.05 100.02 48.65 100.31 ;
      RECT  46.05 28.2 48.65 28.49 ;
      RECT  46.05 89.75 48.65 90.04 ;
      RECT  46.05 53.85 48.65 54.14 ;
      RECT  46.05 64.1 48.65 64.39 ;
      RECT  46.05 74.37 48.65 74.66 ;
      RECT  46.05 64.11 48.65 64.4 ;
      RECT  46.05 94.89 48.65 95.18 ;
      RECT  46.05 43.59 48.65 43.88 ;
      RECT  46.05 105.15 48.65 105.44 ;
      RECT  46.05 84.62 48.65 84.91 ;
      RECT  46.05 84.63 48.65 84.92 ;
      RECT  46.05 33.32 48.65 33.61 ;
      RECT  46.05 53.84 48.65 54.13 ;
      RECT  46.05 43.58 48.65 43.87 ;
      RECT  46.05 105.14 48.65 105.43 ;
      RECT  46.05 74.36 48.65 74.65 ;
      RECT  46.05 115.4 48.65 115.69 ;
      RECT  46.05 33.33 48.65 33.62 ;
      RECT  46.05 94.88 48.65 95.17 ;
      RECT  46.05 15.385 48.65 15.525 ;
      RECT  48.65 15.385 51.25 15.525 ;
      RECT  51.25 15.385 53.85 15.525 ;
      RECT  42.55 15.385 53.85 15.525 ;
      RECT  50.08 8.35 50.37 8.41 ;
      RECT  48.65 8.79 52.65 8.93 ;
      RECT  50.08 8.41 51.54 8.55 ;
      RECT  48.65 12.11 52.65 12.4 ;
      RECT  48.91 9.35 49.22 9.59 ;
      RECT  48.65 10.78 52.65 10.92 ;
      RECT  48.91 9.59 49.2 9.64 ;
      RECT  51.25 8.55 51.54 8.64 ;
      RECT  50.15 9.76 50.48 10.09 ;
      RECT  49.01 10.92 49.3 11.01 ;
      RECT  51.39 9.14 51.72 9.47 ;
      RECT  50.08 8.55 50.37 8.64 ;
      RECT  49.08 8.93 49.22 9.35 ;
      RECT  48.65 7.65 52.65 7.94 ;
      RECT  49.01 10.72 49.3 10.78 ;
      RECT  51.25 8.35 51.54 8.41 ;
      RECT  52.68 8.35 52.97 8.41 ;
      RECT  51.25 8.79 55.25 8.93 ;
      RECT  52.68 8.41 54.14 8.55 ;
      RECT  51.25 12.11 55.25 12.4 ;
      RECT  51.51 9.35 51.82 9.59 ;
      RECT  51.25 10.78 55.25 10.92 ;
      RECT  51.51 9.59 51.8 9.64 ;
      RECT  53.85 8.55 54.14 8.64 ;
      RECT  52.75 9.76 53.08 10.09 ;
      RECT  51.61 10.92 51.9 11.01 ;
      RECT  53.99 9.14 54.32 9.47 ;
      RECT  52.68 8.55 52.97 8.64 ;
      RECT  51.68 8.93 51.82 9.35 ;
      RECT  51.25 7.65 55.25 7.94 ;
      RECT  51.61 10.72 51.9 10.78 ;
      RECT  53.85 8.35 54.14 8.41 ;
      RECT  48.65 10.78 52.65 10.92 ;
      RECT  51.25 10.78 55.25 10.92 ;
      RECT  42.55 9.4 55.25 9.54 ;
      RECT  59.57 4.05 59.87 4.34 ;
      RECT  61.28 1.68 61.58 1.97 ;
      RECT  50.95 2.44 51.25 2.49 ;
      RECT  52.83 2.21 53.12 2.5 ;
      RECT  50.95 2.19 51.25 2.24 ;
      RECT  59.12 2.61 59.45 2.65 ;
      RECT  48.65 1.66 48.95 1.96 ;
      RECT  54.96 3.05 58.79 3.34 ;
      RECT  49.22 2.24 51.25 2.44 ;
      RECT  49.35 -0.17 61.59 0.16 ;
      RECT  53.26 1.72 53.56 4.34 ;
      RECT  59.61 2.01 59.87 4.05 ;
      RECT  49.47 1.68 49.76 1.97 ;
      RECT  54.51 2.32 59.45 2.61 ;
      RECT  61.12 3.05 61.42 3.34 ;
      RECT  59.57 1.72 59.87 2.01 ;
      RECT  49.35 5.58 61.59 6.03 ;
      RECT  62.17 4.05 62.47 4.34 ;
      RECT  63.88 1.68 64.18 1.97 ;
      RECT  53.55 2.44 53.85 2.49 ;
      RECT  55.43 2.21 55.72 2.5 ;
      RECT  53.55 2.19 53.85 2.24 ;
      RECT  61.72 2.61 62.05 2.65 ;
      RECT  51.25 1.66 51.55 1.96 ;
      RECT  57.56 3.05 61.39 3.34 ;
      RECT  51.82 2.24 53.85 2.44 ;
      RECT  51.95 -0.17 64.19 0.16 ;
      RECT  55.86 1.72 56.16 4.34 ;
      RECT  62.21 2.01 62.47 4.05 ;
      RECT  52.07 1.68 52.36 1.97 ;
      RECT  57.11 2.32 62.05 2.61 ;
      RECT  63.72 3.05 64.02 3.34 ;
      RECT  62.17 1.72 62.47 2.01 ;
      RECT  51.95 5.58 64.19 6.03 ;
      RECT  48.65 1.66 48.95 1.96 ;
      RECT  51.25 1.66 51.55 1.96 ;
      RECT  61.28 1.68 61.58 1.97 ;
      RECT  61.12 3.05 61.42 3.34 ;
      RECT  63.88 1.68 64.18 1.97 ;
      RECT  63.72 3.05 64.02 3.34 ;
      RECT  42.55 2.21 64.19 2.35 ;
      RECT  48.65 10.92 52.65 10.78 ;
      RECT  51.25 10.92 55.25 10.78 ;
      RECT  48.65 1.96 48.95 1.66 ;
      RECT  51.25 1.96 51.55 1.66 ;
      RECT  42.55 9.54 55.25 9.4 ;
      RECT  42.55 15.525 53.85 15.385 ;
      RECT  42.55 2.35 64.19 2.21 ;
      RECT  48.65 10.78 52.65 10.92 ;
      RECT  51.25 10.78 55.25 10.92 ;
      RECT  48.65 1.66 48.95 1.96 ;
      RECT  51.25 1.66 51.55 1.96 ;
      RECT  -52.26 -8.84 -47.34 -8.59 ;
      RECT  -55.37 -9.2 -54.69 -8.88 ;
      RECT  -46.46 -8.14 -46.13 -8.02 ;
      RECT  -54.5 -9.32 -54.21 -9.29 ;
      RECT  -55.45 -10.88 -42.92 -10.55 ;
      RECT  -47.54 -9.01 -47.34 -8.84 ;
      RECT  -54.5 -9.09 -54.21 -9.03 ;
      RECT  -46.85 -9.24 -46.55 -9.13 ;
      RECT  -47.54 -8.34 -46.13 -8.14 ;
      RECT  -52.26 -8.35 -51.93 -8.34 ;
      RECT  -48.18 -8.35 -47.85 -8.34 ;
      RECT  -54.22 -8.38 -53.59 -8.06 ;
      RECT  -47.58 -9.34 -47.25 -9.01 ;
      RECT  -53.34 -8.34 -47.85 -8.14 ;
      RECT  -52.65 -9.45 -49.36 -9.24 ;
      RECT  -49.69 -9.5 -49.36 -9.45 ;
      RECT  -48.18 -8.14 -47.85 -8.02 ;
      RECT  -52.26 -8.14 -51.93 -8.02 ;
      RECT  -53.38 -9.09 -53.05 -9.01 ;
      RECT  -52.65 -9.24 -52.35 -9.14 ;
      RECT  -43.66 -9.24 -43.32 -9.21 ;
      RECT  -46.85 -9.44 -43.32 -9.24 ;
      RECT  -49.69 -9.24 -49.36 -9.17 ;
      RECT  -45.32 -8.69 -44.69 -8.37 ;
      RECT  -52.26 -8.59 -51.93 -8.56 ;
      RECT  -53.38 -9.34 -53.05 -9.29 ;
      RECT  -43.66 -9.54 -43.32 -9.44 ;
      RECT  -46.46 -8.35 -46.13 -8.34 ;
      RECT  -52.26 -8.89 -51.93 -8.84 ;
      RECT  -54.5 -9.29 -53.05 -9.09 ;
      RECT  -55.39 -6.79 -42.74 -6.46 ;
      RECT  -53.34 -9.01 -53.14 -8.34 ;
      RECT  -47.54 -8.59 -47.34 -8.34 ;
      RECT  -55.39 -6.79 -31.52 -6.46 ;
      RECT  -55.45 -10.88 -31.58 -10.55 ;
      RECT  -52.26 -4.4 -47.34 -4.65 ;
      RECT  -55.37 -4.04 -54.69 -4.36 ;
      RECT  -46.46 -5.1 -46.13 -5.22 ;
      RECT  -54.5 -3.92 -54.21 -3.95 ;
      RECT  -55.45 -2.36 -42.92 -2.69 ;
      RECT  -47.54 -4.23 -47.34 -4.4 ;
      RECT  -54.5 -4.15 -54.21 -4.21 ;
      RECT  -46.85 -4.0 -46.55 -4.11 ;
      RECT  -47.54 -4.9 -46.13 -5.1 ;
      RECT  -52.26 -4.89 -51.93 -4.9 ;
      RECT  -48.18 -4.89 -47.85 -4.9 ;
      RECT  -54.22 -4.86 -53.59 -5.18 ;
      RECT  -47.58 -3.9 -47.25 -4.23 ;
      RECT  -53.34 -4.9 -47.85 -5.1 ;
      RECT  -52.65 -3.79 -49.36 -4.0 ;
      RECT  -49.69 -3.74 -49.36 -3.79 ;
      RECT  -48.18 -5.1 -47.85 -5.22 ;
      RECT  -52.26 -5.1 -51.93 -5.22 ;
      RECT  -53.38 -4.15 -53.05 -4.23 ;
      RECT  -52.65 -4.0 -52.35 -4.1 ;
      RECT  -43.66 -4.0 -43.32 -4.03 ;
      RECT  -46.85 -3.8 -43.32 -4.0 ;
      RECT  -49.69 -4.0 -49.36 -4.07 ;
      RECT  -45.32 -4.55 -44.69 -4.87 ;
      RECT  -52.26 -4.65 -51.93 -4.68 ;
      RECT  -53.38 -3.9 -53.05 -3.95 ;
      RECT  -43.66 -3.7 -43.32 -3.8 ;
      RECT  -46.46 -4.89 -46.13 -4.9 ;
      RECT  -52.26 -4.35 -51.93 -4.4 ;
      RECT  -54.5 -3.95 -53.05 -4.15 ;
      RECT  -55.39 -6.45 -42.74 -6.78 ;
      RECT  -53.34 -4.23 -53.14 -4.9 ;
      RECT  -47.54 -4.65 -47.34 -4.9 ;
      RECT  -55.39 -6.45 -31.52 -6.78 ;
      RECT  -55.45 -2.36 -31.58 -2.69 ;
      RECT  -10.84 101.88 -5.92 102.13 ;
      RECT  -13.95 101.52 -13.27 101.84 ;
      RECT  -5.04 102.58 -4.71 102.7 ;
      RECT  -13.08 101.4 -12.79 101.43 ;
      RECT  -14.03 99.84 -1.5 100.17 ;
      RECT  -6.12 101.71 -5.92 101.88 ;
      RECT  -13.08 101.63 -12.79 101.69 ;
      RECT  -5.43 101.48 -5.13 101.59 ;
      RECT  -6.12 102.38 -4.71 102.58 ;
      RECT  -10.84 102.37 -10.51 102.38 ;
      RECT  -6.76 102.37 -6.43 102.38 ;
      RECT  -12.8 102.34 -12.17 102.66 ;
      RECT  -6.16 101.38 -5.83 101.71 ;
      RECT  -11.92 102.38 -6.43 102.58 ;
      RECT  -11.23 101.27 -7.94 101.48 ;
      RECT  -8.27 101.22 -7.94 101.27 ;
      RECT  -6.76 102.58 -6.43 102.7 ;
      RECT  -10.84 102.58 -10.51 102.7 ;
      RECT  -11.96 101.63 -11.63 101.71 ;
      RECT  -11.23 101.48 -10.93 101.58 ;
      RECT  -2.24 101.48 -1.9 101.51 ;
      RECT  -5.43 101.28 -1.9 101.48 ;
      RECT  -8.27 101.48 -7.94 101.55 ;
      RECT  -3.9 102.03 -3.27 102.35 ;
      RECT  -10.84 102.13 -10.51 102.16 ;
      RECT  -11.96 101.38 -11.63 101.43 ;
      RECT  -2.24 101.18 -1.9 101.28 ;
      RECT  -5.04 102.37 -4.71 102.38 ;
      RECT  -10.84 101.83 -10.51 101.88 ;
      RECT  -13.08 101.43 -11.63 101.63 ;
      RECT  -13.97 103.93 -1.32 104.26 ;
      RECT  -11.92 101.71 -11.72 102.38 ;
      RECT  -6.12 102.13 -5.92 102.38 ;
      RECT  -10.84 106.32 -5.92 106.07 ;
      RECT  -13.95 106.68 -13.27 106.36 ;
      RECT  -5.04 105.62 -4.71 105.5 ;
      RECT  -13.08 106.8 -12.79 106.77 ;
      RECT  -14.03 108.36 -1.5 108.03 ;
      RECT  -6.12 106.49 -5.92 106.32 ;
      RECT  -13.08 106.57 -12.79 106.51 ;
      RECT  -5.43 106.72 -5.13 106.61 ;
      RECT  -6.12 105.82 -4.71 105.62 ;
      RECT  -10.84 105.83 -10.51 105.82 ;
      RECT  -6.76 105.83 -6.43 105.82 ;
      RECT  -12.8 105.86 -12.17 105.54 ;
      RECT  -6.16 106.82 -5.83 106.49 ;
      RECT  -11.92 105.82 -6.43 105.62 ;
      RECT  -11.23 106.93 -7.94 106.72 ;
      RECT  -8.27 106.98 -7.94 106.93 ;
      RECT  -6.76 105.62 -6.43 105.5 ;
      RECT  -10.84 105.62 -10.51 105.5 ;
      RECT  -11.96 106.57 -11.63 106.49 ;
      RECT  -11.23 106.72 -10.93 106.62 ;
      RECT  -2.24 106.72 -1.9 106.69 ;
      RECT  -5.43 106.92 -1.9 106.72 ;
      RECT  -8.27 106.72 -7.94 106.65 ;
      RECT  -3.9 106.17 -3.27 105.85 ;
      RECT  -10.84 106.07 -10.51 106.04 ;
      RECT  -11.96 106.82 -11.63 106.77 ;
      RECT  -2.24 107.02 -1.9 106.92 ;
      RECT  -5.04 105.83 -4.71 105.82 ;
      RECT  -10.84 106.37 -10.51 106.32 ;
      RECT  -13.08 106.77 -11.63 106.57 ;
      RECT  -13.97 104.27 -1.32 103.94 ;
      RECT  -11.92 106.49 -11.72 105.82 ;
      RECT  -6.12 106.07 -5.92 105.82 ;
      RECT  -10.84 110.06 -5.92 110.31 ;
      RECT  -13.95 109.7 -13.27 110.02 ;
      RECT  -5.04 110.76 -4.71 110.88 ;
      RECT  -13.08 109.58 -12.79 109.61 ;
      RECT  -14.03 108.02 -1.5 108.35 ;
      RECT  -6.12 109.89 -5.92 110.06 ;
      RECT  -13.08 109.81 -12.79 109.87 ;
      RECT  -5.43 109.66 -5.13 109.77 ;
      RECT  -6.12 110.56 -4.71 110.76 ;
      RECT  -10.84 110.55 -10.51 110.56 ;
      RECT  -6.76 110.55 -6.43 110.56 ;
      RECT  -12.8 110.52 -12.17 110.84 ;
      RECT  -6.16 109.56 -5.83 109.89 ;
      RECT  -11.92 110.56 -6.43 110.76 ;
      RECT  -11.23 109.45 -7.94 109.66 ;
      RECT  -8.27 109.4 -7.94 109.45 ;
      RECT  -6.76 110.76 -6.43 110.88 ;
      RECT  -10.84 110.76 -10.51 110.88 ;
      RECT  -11.96 109.81 -11.63 109.89 ;
      RECT  -11.23 109.66 -10.93 109.76 ;
      RECT  -2.24 109.66 -1.9 109.69 ;
      RECT  -5.43 109.46 -1.9 109.66 ;
      RECT  -8.27 109.66 -7.94 109.73 ;
      RECT  -3.9 110.21 -3.27 110.53 ;
      RECT  -10.84 110.31 -10.51 110.34 ;
      RECT  -11.96 109.56 -11.63 109.61 ;
      RECT  -2.24 109.36 -1.9 109.46 ;
      RECT  -5.04 110.55 -4.71 110.56 ;
      RECT  -10.84 110.01 -10.51 110.06 ;
      RECT  -13.08 109.61 -11.63 109.81 ;
      RECT  -13.97 112.11 -1.32 112.44 ;
      RECT  -11.92 109.89 -11.72 110.56 ;
      RECT  -6.12 110.31 -5.92 110.56 ;
      RECT  -10.84 114.5 -5.92 114.25 ;
      RECT  -13.95 114.86 -13.27 114.54 ;
      RECT  -5.04 113.8 -4.71 113.68 ;
      RECT  -13.08 114.98 -12.79 114.95 ;
      RECT  -14.03 116.54 -1.5 116.21 ;
      RECT  -6.12 114.67 -5.92 114.5 ;
      RECT  -13.08 114.75 -12.79 114.69 ;
      RECT  -5.43 114.9 -5.13 114.79 ;
      RECT  -6.12 114.0 -4.71 113.8 ;
      RECT  -10.84 114.01 -10.51 114.0 ;
      RECT  -6.76 114.01 -6.43 114.0 ;
      RECT  -12.8 114.04 -12.17 113.72 ;
      RECT  -6.16 115.0 -5.83 114.67 ;
      RECT  -11.92 114.0 -6.43 113.8 ;
      RECT  -11.23 115.11 -7.94 114.9 ;
      RECT  -8.27 115.16 -7.94 115.11 ;
      RECT  -6.76 113.8 -6.43 113.68 ;
      RECT  -10.84 113.8 -10.51 113.68 ;
      RECT  -11.96 114.75 -11.63 114.67 ;
      RECT  -11.23 114.9 -10.93 114.8 ;
      RECT  -2.24 114.9 -1.9 114.87 ;
      RECT  -5.43 115.1 -1.9 114.9 ;
      RECT  -8.27 114.9 -7.94 114.83 ;
      RECT  -3.9 114.35 -3.27 114.03 ;
      RECT  -10.84 114.25 -10.51 114.22 ;
      RECT  -11.96 115.0 -11.63 114.95 ;
      RECT  -2.24 115.2 -1.9 115.1 ;
      RECT  -5.04 114.01 -4.71 114.0 ;
      RECT  -10.84 114.55 -10.51 114.5 ;
      RECT  -13.08 114.95 -11.63 114.75 ;
      RECT  -13.97 112.45 -1.32 112.12 ;
      RECT  -11.92 114.67 -11.72 114.0 ;
      RECT  -6.12 114.25 -5.92 114.0 ;
      RECT  14.58 -8.84 19.5 -8.59 ;
      RECT  11.47 -9.2 12.15 -8.88 ;
      RECT  20.38 -8.14 20.71 -8.02 ;
      RECT  12.34 -9.32 12.63 -9.29 ;
      RECT  11.39 -10.88 23.92 -10.55 ;
      RECT  19.3 -9.01 19.5 -8.84 ;
      RECT  12.34 -9.09 12.63 -9.03 ;
      RECT  19.99 -9.24 20.29 -9.13 ;
      RECT  19.3 -8.34 20.71 -8.14 ;
      RECT  14.58 -8.35 14.91 -8.34 ;
      RECT  18.66 -8.35 18.99 -8.34 ;
      RECT  12.62 -8.38 13.25 -8.06 ;
      RECT  19.26 -9.34 19.59 -9.01 ;
      RECT  13.5 -8.34 18.99 -8.14 ;
      RECT  14.19 -9.45 17.48 -9.24 ;
      RECT  17.15 -9.5 17.48 -9.45 ;
      RECT  18.66 -8.14 18.99 -8.02 ;
      RECT  14.58 -8.14 14.91 -8.02 ;
      RECT  13.46 -9.09 13.79 -9.01 ;
      RECT  14.19 -9.24 14.49 -9.14 ;
      RECT  23.18 -9.24 23.52 -9.21 ;
      RECT  19.99 -9.44 23.52 -9.24 ;
      RECT  17.15 -9.24 17.48 -9.17 ;
      RECT  21.52 -8.69 22.15 -8.37 ;
      RECT  14.58 -8.59 14.91 -8.56 ;
      RECT  13.46 -9.34 13.79 -9.29 ;
      RECT  23.18 -9.54 23.52 -9.44 ;
      RECT  20.38 -8.35 20.71 -8.34 ;
      RECT  14.58 -8.89 14.91 -8.84 ;
      RECT  12.34 -9.29 13.79 -9.09 ;
      RECT  11.45 -6.79 24.1 -6.46 ;
      RECT  13.5 -9.01 13.7 -8.34 ;
      RECT  19.3 -8.59 19.5 -8.34 ;
      RECT  27.29 -8.84 32.21 -8.59 ;
      RECT  24.18 -9.2 24.86 -8.88 ;
      RECT  33.09 -8.14 33.42 -8.02 ;
      RECT  25.05 -9.32 25.34 -9.29 ;
      RECT  24.1 -10.88 36.63 -10.55 ;
      RECT  32.01 -9.01 32.21 -8.84 ;
      RECT  25.05 -9.09 25.34 -9.03 ;
      RECT  32.7 -9.24 33.0 -9.13 ;
      RECT  32.01 -8.34 33.42 -8.14 ;
      RECT  27.29 -8.35 27.62 -8.34 ;
      RECT  31.37 -8.35 31.7 -8.34 ;
      RECT  25.33 -8.38 25.96 -8.06 ;
      RECT  31.97 -9.34 32.3 -9.01 ;
      RECT  26.21 -8.34 31.7 -8.14 ;
      RECT  26.9 -9.45 30.19 -9.24 ;
      RECT  29.86 -9.5 30.19 -9.45 ;
      RECT  31.37 -8.14 31.7 -8.02 ;
      RECT  27.29 -8.14 27.62 -8.02 ;
      RECT  26.17 -9.09 26.5 -9.01 ;
      RECT  26.9 -9.24 27.2 -9.14 ;
      RECT  35.89 -9.24 36.23 -9.21 ;
      RECT  32.7 -9.44 36.23 -9.24 ;
      RECT  29.86 -9.24 30.19 -9.17 ;
      RECT  34.23 -8.69 34.86 -8.37 ;
      RECT  27.29 -8.59 27.62 -8.56 ;
      RECT  26.17 -9.34 26.5 -9.29 ;
      RECT  35.89 -9.54 36.23 -9.44 ;
      RECT  33.09 -8.35 33.42 -8.34 ;
      RECT  27.29 -8.89 27.62 -8.84 ;
      RECT  25.05 -9.29 26.5 -9.09 ;
      RECT  24.16 -6.79 36.81 -6.46 ;
      RECT  26.21 -9.01 26.41 -8.34 ;
      RECT  32.01 -8.59 32.21 -8.34 ;
   LAYER  m2 ;
      RECT  50.49 34.17 50.63 39.07 ;
      RECT  49.78 33.26 50.21 33.69 ;
      RECT  49.37 34.17 49.51 39.05 ;
      RECT  50.49 33.82 50.84 34.17 ;
      RECT  49.16 33.82 49.51 34.17 ;
      RECT  49.37 33.17 49.51 33.82 ;
      RECT  50.49 33.17 50.63 33.82 ;
      RECT  49.78 38.38 50.21 38.81 ;
      RECT  50.49 43.03 50.63 38.13 ;
      RECT  49.78 43.94 50.21 43.51 ;
      RECT  49.37 43.03 49.51 38.15 ;
      RECT  50.49 43.38 50.84 43.03 ;
      RECT  49.16 43.38 49.51 43.03 ;
      RECT  49.37 44.03 49.51 43.38 ;
      RECT  50.49 44.03 50.63 43.38 ;
      RECT  49.78 38.82 50.21 38.39 ;
      RECT  50.49 44.43 50.63 49.33 ;
      RECT  49.78 43.52 50.21 43.95 ;
      RECT  49.37 44.43 49.51 49.31 ;
      RECT  50.49 44.08 50.84 44.43 ;
      RECT  49.16 44.08 49.51 44.43 ;
      RECT  49.37 43.43 49.51 44.08 ;
      RECT  50.49 43.43 50.63 44.08 ;
      RECT  49.78 48.64 50.21 49.07 ;
      RECT  50.49 53.29 50.63 48.39 ;
      RECT  49.78 54.2 50.21 53.77 ;
      RECT  49.37 53.29 49.51 48.41 ;
      RECT  50.49 53.64 50.84 53.29 ;
      RECT  49.16 53.64 49.51 53.29 ;
      RECT  49.37 54.29 49.51 53.64 ;
      RECT  50.49 54.29 50.63 53.64 ;
      RECT  49.78 49.08 50.21 48.65 ;
      RECT  50.49 54.69 50.63 59.59 ;
      RECT  49.78 53.78 50.21 54.21 ;
      RECT  49.37 54.69 49.51 59.57 ;
      RECT  50.49 54.34 50.84 54.69 ;
      RECT  49.16 54.34 49.51 54.69 ;
      RECT  49.37 53.69 49.51 54.34 ;
      RECT  50.49 53.69 50.63 54.34 ;
      RECT  49.78 58.9 50.21 59.33 ;
      RECT  50.49 63.55 50.63 58.65 ;
      RECT  49.78 64.46 50.21 64.03 ;
      RECT  49.37 63.55 49.51 58.67 ;
      RECT  50.49 63.9 50.84 63.55 ;
      RECT  49.16 63.9 49.51 63.55 ;
      RECT  49.37 64.55 49.51 63.9 ;
      RECT  50.49 64.55 50.63 63.9 ;
      RECT  49.78 59.34 50.21 58.91 ;
      RECT  50.49 64.95 50.63 69.85 ;
      RECT  49.78 64.04 50.21 64.47 ;
      RECT  49.37 64.95 49.51 69.83 ;
      RECT  50.49 64.6 50.84 64.95 ;
      RECT  49.16 64.6 49.51 64.95 ;
      RECT  49.37 63.95 49.51 64.6 ;
      RECT  50.49 63.95 50.63 64.6 ;
      RECT  49.78 69.16 50.21 69.59 ;
      RECT  50.49 73.81 50.63 68.91 ;
      RECT  49.78 74.72 50.21 74.29 ;
      RECT  49.37 73.81 49.51 68.93 ;
      RECT  50.49 74.16 50.84 73.81 ;
      RECT  49.16 74.16 49.51 73.81 ;
      RECT  49.37 74.81 49.51 74.16 ;
      RECT  50.49 74.81 50.63 74.16 ;
      RECT  49.78 69.6 50.21 69.17 ;
      RECT  50.49 75.21 50.63 80.11 ;
      RECT  49.78 74.3 50.21 74.73 ;
      RECT  49.37 75.21 49.51 80.09 ;
      RECT  50.49 74.86 50.84 75.21 ;
      RECT  49.16 74.86 49.51 75.21 ;
      RECT  49.37 74.21 49.51 74.86 ;
      RECT  50.49 74.21 50.63 74.86 ;
      RECT  49.78 79.42 50.21 79.85 ;
      RECT  50.49 84.07 50.63 79.17 ;
      RECT  49.78 84.98 50.21 84.55 ;
      RECT  49.37 84.07 49.51 79.19 ;
      RECT  50.49 84.42 50.84 84.07 ;
      RECT  49.16 84.42 49.51 84.07 ;
      RECT  49.37 85.07 49.51 84.42 ;
      RECT  50.49 85.07 50.63 84.42 ;
      RECT  49.78 79.86 50.21 79.43 ;
      RECT  50.49 85.47 50.63 90.37 ;
      RECT  49.78 84.56 50.21 84.99 ;
      RECT  49.37 85.47 49.51 90.35 ;
      RECT  50.49 85.12 50.84 85.47 ;
      RECT  49.16 85.12 49.51 85.47 ;
      RECT  49.37 84.47 49.51 85.12 ;
      RECT  50.49 84.47 50.63 85.12 ;
      RECT  49.78 89.68 50.21 90.11 ;
      RECT  50.49 94.33 50.63 89.43 ;
      RECT  49.78 95.24 50.21 94.81 ;
      RECT  49.37 94.33 49.51 89.45 ;
      RECT  50.49 94.68 50.84 94.33 ;
      RECT  49.16 94.68 49.51 94.33 ;
      RECT  49.37 95.33 49.51 94.68 ;
      RECT  50.49 95.33 50.63 94.68 ;
      RECT  49.78 90.12 50.21 89.69 ;
      RECT  50.49 95.73 50.63 100.63 ;
      RECT  49.78 94.82 50.21 95.25 ;
      RECT  49.37 95.73 49.51 100.61 ;
      RECT  50.49 95.38 50.84 95.73 ;
      RECT  49.16 95.38 49.51 95.73 ;
      RECT  49.37 94.73 49.51 95.38 ;
      RECT  50.49 94.73 50.63 95.38 ;
      RECT  49.78 99.94 50.21 100.37 ;
      RECT  50.49 104.59 50.63 99.69 ;
      RECT  49.78 105.5 50.21 105.07 ;
      RECT  49.37 104.59 49.51 99.71 ;
      RECT  50.49 104.94 50.84 104.59 ;
      RECT  49.16 104.94 49.51 104.59 ;
      RECT  49.37 105.59 49.51 104.94 ;
      RECT  50.49 105.59 50.63 104.94 ;
      RECT  49.78 100.38 50.21 99.95 ;
      RECT  50.49 105.99 50.63 110.89 ;
      RECT  49.78 105.08 50.21 105.51 ;
      RECT  49.37 105.99 49.51 110.87 ;
      RECT  50.49 105.64 50.84 105.99 ;
      RECT  49.16 105.64 49.51 105.99 ;
      RECT  49.37 104.99 49.51 105.64 ;
      RECT  50.49 104.99 50.63 105.64 ;
      RECT  49.78 110.2 50.21 110.63 ;
      RECT  50.49 114.85 50.63 109.95 ;
      RECT  49.78 115.76 50.21 115.33 ;
      RECT  49.37 114.85 49.51 109.97 ;
      RECT  50.49 115.2 50.84 114.85 ;
      RECT  49.16 115.2 49.51 114.85 ;
      RECT  49.37 115.85 49.51 115.2 ;
      RECT  50.49 115.85 50.63 115.2 ;
      RECT  49.78 110.64 50.21 110.21 ;
      RECT  53.09 34.17 53.23 39.07 ;
      RECT  52.38 33.26 52.81 33.69 ;
      RECT  51.97 34.17 52.11 39.05 ;
      RECT  53.09 33.82 53.44 34.17 ;
      RECT  51.76 33.82 52.11 34.17 ;
      RECT  51.97 33.17 52.11 33.82 ;
      RECT  53.09 33.17 53.23 33.82 ;
      RECT  52.38 38.38 52.81 38.81 ;
      RECT  53.09 43.03 53.23 38.13 ;
      RECT  52.38 43.94 52.81 43.51 ;
      RECT  51.97 43.03 52.11 38.15 ;
      RECT  53.09 43.38 53.44 43.03 ;
      RECT  51.76 43.38 52.11 43.03 ;
      RECT  51.97 44.03 52.11 43.38 ;
      RECT  53.09 44.03 53.23 43.38 ;
      RECT  52.38 38.82 52.81 38.39 ;
      RECT  53.09 44.43 53.23 49.33 ;
      RECT  52.38 43.52 52.81 43.95 ;
      RECT  51.97 44.43 52.11 49.31 ;
      RECT  53.09 44.08 53.44 44.43 ;
      RECT  51.76 44.08 52.11 44.43 ;
      RECT  51.97 43.43 52.11 44.08 ;
      RECT  53.09 43.43 53.23 44.08 ;
      RECT  52.38 48.64 52.81 49.07 ;
      RECT  53.09 53.29 53.23 48.39 ;
      RECT  52.38 54.2 52.81 53.77 ;
      RECT  51.97 53.29 52.11 48.41 ;
      RECT  53.09 53.64 53.44 53.29 ;
      RECT  51.76 53.64 52.11 53.29 ;
      RECT  51.97 54.29 52.11 53.64 ;
      RECT  53.09 54.29 53.23 53.64 ;
      RECT  52.38 49.08 52.81 48.65 ;
      RECT  53.09 54.69 53.23 59.59 ;
      RECT  52.38 53.78 52.81 54.21 ;
      RECT  51.97 54.69 52.11 59.57 ;
      RECT  53.09 54.34 53.44 54.69 ;
      RECT  51.76 54.34 52.11 54.69 ;
      RECT  51.97 53.69 52.11 54.34 ;
      RECT  53.09 53.69 53.23 54.34 ;
      RECT  52.38 58.9 52.81 59.33 ;
      RECT  53.09 63.55 53.23 58.65 ;
      RECT  52.38 64.46 52.81 64.03 ;
      RECT  51.97 63.55 52.11 58.67 ;
      RECT  53.09 63.9 53.44 63.55 ;
      RECT  51.76 63.9 52.11 63.55 ;
      RECT  51.97 64.55 52.11 63.9 ;
      RECT  53.09 64.55 53.23 63.9 ;
      RECT  52.38 59.34 52.81 58.91 ;
      RECT  53.09 64.95 53.23 69.85 ;
      RECT  52.38 64.04 52.81 64.47 ;
      RECT  51.97 64.95 52.11 69.83 ;
      RECT  53.09 64.6 53.44 64.95 ;
      RECT  51.76 64.6 52.11 64.95 ;
      RECT  51.97 63.95 52.11 64.6 ;
      RECT  53.09 63.95 53.23 64.6 ;
      RECT  52.38 69.16 52.81 69.59 ;
      RECT  53.09 73.81 53.23 68.91 ;
      RECT  52.38 74.72 52.81 74.29 ;
      RECT  51.97 73.81 52.11 68.93 ;
      RECT  53.09 74.16 53.44 73.81 ;
      RECT  51.76 74.16 52.11 73.81 ;
      RECT  51.97 74.81 52.11 74.16 ;
      RECT  53.09 74.81 53.23 74.16 ;
      RECT  52.38 69.6 52.81 69.17 ;
      RECT  53.09 75.21 53.23 80.11 ;
      RECT  52.38 74.3 52.81 74.73 ;
      RECT  51.97 75.21 52.11 80.09 ;
      RECT  53.09 74.86 53.44 75.21 ;
      RECT  51.76 74.86 52.11 75.21 ;
      RECT  51.97 74.21 52.11 74.86 ;
      RECT  53.09 74.21 53.23 74.86 ;
      RECT  52.38 79.42 52.81 79.85 ;
      RECT  53.09 84.07 53.23 79.17 ;
      RECT  52.38 84.98 52.81 84.55 ;
      RECT  51.97 84.07 52.11 79.19 ;
      RECT  53.09 84.42 53.44 84.07 ;
      RECT  51.76 84.42 52.11 84.07 ;
      RECT  51.97 85.07 52.11 84.42 ;
      RECT  53.09 85.07 53.23 84.42 ;
      RECT  52.38 79.86 52.81 79.43 ;
      RECT  53.09 85.47 53.23 90.37 ;
      RECT  52.38 84.56 52.81 84.99 ;
      RECT  51.97 85.47 52.11 90.35 ;
      RECT  53.09 85.12 53.44 85.47 ;
      RECT  51.76 85.12 52.11 85.47 ;
      RECT  51.97 84.47 52.11 85.12 ;
      RECT  53.09 84.47 53.23 85.12 ;
      RECT  52.38 89.68 52.81 90.11 ;
      RECT  53.09 94.33 53.23 89.43 ;
      RECT  52.38 95.24 52.81 94.81 ;
      RECT  51.97 94.33 52.11 89.45 ;
      RECT  53.09 94.68 53.44 94.33 ;
      RECT  51.76 94.68 52.11 94.33 ;
      RECT  51.97 95.33 52.11 94.68 ;
      RECT  53.09 95.33 53.23 94.68 ;
      RECT  52.38 90.12 52.81 89.69 ;
      RECT  53.09 95.73 53.23 100.63 ;
      RECT  52.38 94.82 52.81 95.25 ;
      RECT  51.97 95.73 52.11 100.61 ;
      RECT  53.09 95.38 53.44 95.73 ;
      RECT  51.76 95.38 52.11 95.73 ;
      RECT  51.97 94.73 52.11 95.38 ;
      RECT  53.09 94.73 53.23 95.38 ;
      RECT  52.38 99.94 52.81 100.37 ;
      RECT  53.09 104.59 53.23 99.69 ;
      RECT  52.38 105.5 52.81 105.07 ;
      RECT  51.97 104.59 52.11 99.71 ;
      RECT  53.09 104.94 53.44 104.59 ;
      RECT  51.76 104.94 52.11 104.59 ;
      RECT  51.97 105.59 52.11 104.94 ;
      RECT  53.09 105.59 53.23 104.94 ;
      RECT  52.38 100.38 52.81 99.95 ;
      RECT  53.09 105.99 53.23 110.89 ;
      RECT  52.38 105.08 52.81 105.51 ;
      RECT  51.97 105.99 52.11 110.87 ;
      RECT  53.09 105.64 53.44 105.99 ;
      RECT  51.76 105.64 52.11 105.99 ;
      RECT  51.97 104.99 52.11 105.64 ;
      RECT  53.09 104.99 53.23 105.64 ;
      RECT  52.38 110.2 52.81 110.63 ;
      RECT  53.09 114.85 53.23 109.95 ;
      RECT  52.38 115.76 52.81 115.33 ;
      RECT  51.97 114.85 52.11 109.97 ;
      RECT  53.09 115.2 53.44 114.85 ;
      RECT  51.76 115.2 52.11 114.85 ;
      RECT  51.97 115.85 52.11 115.2 ;
      RECT  53.09 115.85 53.23 115.2 ;
      RECT  52.38 110.64 52.81 110.21 ;
      RECT  49.37 33.47 49.51 115.55 ;
      RECT  50.49 33.47 50.63 115.55 ;
      RECT  51.97 33.47 52.11 115.55 ;
      RECT  53.09 33.47 53.23 115.55 ;
      RECT  47.89 23.91 48.03 28.81 ;
      RECT  47.18 23.0 47.61 23.43 ;
      RECT  46.77 23.91 46.91 28.79 ;
      RECT  47.89 23.56 48.24 23.91 ;
      RECT  46.56 23.56 46.91 23.91 ;
      RECT  46.77 22.91 46.91 23.56 ;
      RECT  47.89 22.91 48.03 23.56 ;
      RECT  47.18 28.12 47.61 28.55 ;
      RECT  47.89 32.77 48.03 27.87 ;
      RECT  47.18 33.68 47.61 33.25 ;
      RECT  46.77 32.77 46.91 27.89 ;
      RECT  47.89 33.12 48.24 32.77 ;
      RECT  46.56 33.12 46.91 32.77 ;
      RECT  46.77 33.77 46.91 33.12 ;
      RECT  47.89 33.77 48.03 33.12 ;
      RECT  47.18 28.56 47.61 28.13 ;
      RECT  47.89 34.17 48.03 39.07 ;
      RECT  47.18 33.26 47.61 33.69 ;
      RECT  46.77 34.17 46.91 39.05 ;
      RECT  47.89 33.82 48.24 34.17 ;
      RECT  46.56 33.82 46.91 34.17 ;
      RECT  46.77 33.17 46.91 33.82 ;
      RECT  47.89 33.17 48.03 33.82 ;
      RECT  47.18 38.38 47.61 38.81 ;
      RECT  47.89 43.03 48.03 38.13 ;
      RECT  47.18 43.94 47.61 43.51 ;
      RECT  46.77 43.03 46.91 38.15 ;
      RECT  47.89 43.38 48.24 43.03 ;
      RECT  46.56 43.38 46.91 43.03 ;
      RECT  46.77 44.03 46.91 43.38 ;
      RECT  47.89 44.03 48.03 43.38 ;
      RECT  47.18 38.82 47.61 38.39 ;
      RECT  47.89 44.43 48.03 49.33 ;
      RECT  47.18 43.52 47.61 43.95 ;
      RECT  46.77 44.43 46.91 49.31 ;
      RECT  47.89 44.08 48.24 44.43 ;
      RECT  46.56 44.08 46.91 44.43 ;
      RECT  46.77 43.43 46.91 44.08 ;
      RECT  47.89 43.43 48.03 44.08 ;
      RECT  47.18 48.64 47.61 49.07 ;
      RECT  47.89 53.29 48.03 48.39 ;
      RECT  47.18 54.2 47.61 53.77 ;
      RECT  46.77 53.29 46.91 48.41 ;
      RECT  47.89 53.64 48.24 53.29 ;
      RECT  46.56 53.64 46.91 53.29 ;
      RECT  46.77 54.29 46.91 53.64 ;
      RECT  47.89 54.29 48.03 53.64 ;
      RECT  47.18 49.08 47.61 48.65 ;
      RECT  47.89 54.69 48.03 59.59 ;
      RECT  47.18 53.78 47.61 54.21 ;
      RECT  46.77 54.69 46.91 59.57 ;
      RECT  47.89 54.34 48.24 54.69 ;
      RECT  46.56 54.34 46.91 54.69 ;
      RECT  46.77 53.69 46.91 54.34 ;
      RECT  47.89 53.69 48.03 54.34 ;
      RECT  47.18 58.9 47.61 59.33 ;
      RECT  47.89 63.55 48.03 58.65 ;
      RECT  47.18 64.46 47.61 64.03 ;
      RECT  46.77 63.55 46.91 58.67 ;
      RECT  47.89 63.9 48.24 63.55 ;
      RECT  46.56 63.9 46.91 63.55 ;
      RECT  46.77 64.55 46.91 63.9 ;
      RECT  47.89 64.55 48.03 63.9 ;
      RECT  47.18 59.34 47.61 58.91 ;
      RECT  47.89 64.95 48.03 69.85 ;
      RECT  47.18 64.04 47.61 64.47 ;
      RECT  46.77 64.95 46.91 69.83 ;
      RECT  47.89 64.6 48.24 64.95 ;
      RECT  46.56 64.6 46.91 64.95 ;
      RECT  46.77 63.95 46.91 64.6 ;
      RECT  47.89 63.95 48.03 64.6 ;
      RECT  47.18 69.16 47.61 69.59 ;
      RECT  47.89 73.81 48.03 68.91 ;
      RECT  47.18 74.72 47.61 74.29 ;
      RECT  46.77 73.81 46.91 68.93 ;
      RECT  47.89 74.16 48.24 73.81 ;
      RECT  46.56 74.16 46.91 73.81 ;
      RECT  46.77 74.81 46.91 74.16 ;
      RECT  47.89 74.81 48.03 74.16 ;
      RECT  47.18 69.6 47.61 69.17 ;
      RECT  47.89 75.21 48.03 80.11 ;
      RECT  47.18 74.3 47.61 74.73 ;
      RECT  46.77 75.21 46.91 80.09 ;
      RECT  47.89 74.86 48.24 75.21 ;
      RECT  46.56 74.86 46.91 75.21 ;
      RECT  46.77 74.21 46.91 74.86 ;
      RECT  47.89 74.21 48.03 74.86 ;
      RECT  47.18 79.42 47.61 79.85 ;
      RECT  47.89 84.07 48.03 79.17 ;
      RECT  47.18 84.98 47.61 84.55 ;
      RECT  46.77 84.07 46.91 79.19 ;
      RECT  47.89 84.42 48.24 84.07 ;
      RECT  46.56 84.42 46.91 84.07 ;
      RECT  46.77 85.07 46.91 84.42 ;
      RECT  47.89 85.07 48.03 84.42 ;
      RECT  47.18 79.86 47.61 79.43 ;
      RECT  47.89 85.47 48.03 90.37 ;
      RECT  47.18 84.56 47.61 84.99 ;
      RECT  46.77 85.47 46.91 90.35 ;
      RECT  47.89 85.12 48.24 85.47 ;
      RECT  46.56 85.12 46.91 85.47 ;
      RECT  46.77 84.47 46.91 85.12 ;
      RECT  47.89 84.47 48.03 85.12 ;
      RECT  47.18 89.68 47.61 90.11 ;
      RECT  47.89 94.33 48.03 89.43 ;
      RECT  47.18 95.24 47.61 94.81 ;
      RECT  46.77 94.33 46.91 89.45 ;
      RECT  47.89 94.68 48.24 94.33 ;
      RECT  46.56 94.68 46.91 94.33 ;
      RECT  46.77 95.33 46.91 94.68 ;
      RECT  47.89 95.33 48.03 94.68 ;
      RECT  47.18 90.12 47.61 89.69 ;
      RECT  47.89 95.73 48.03 100.63 ;
      RECT  47.18 94.82 47.61 95.25 ;
      RECT  46.77 95.73 46.91 100.61 ;
      RECT  47.89 95.38 48.24 95.73 ;
      RECT  46.56 95.38 46.91 95.73 ;
      RECT  46.77 94.73 46.91 95.38 ;
      RECT  47.89 94.73 48.03 95.38 ;
      RECT  47.18 99.94 47.61 100.37 ;
      RECT  47.89 104.59 48.03 99.69 ;
      RECT  47.18 105.5 47.61 105.07 ;
      RECT  46.77 104.59 46.91 99.71 ;
      RECT  47.89 104.94 48.24 104.59 ;
      RECT  46.56 104.94 46.91 104.59 ;
      RECT  46.77 105.59 46.91 104.94 ;
      RECT  47.89 105.59 48.03 104.94 ;
      RECT  47.18 100.38 47.61 99.95 ;
      RECT  47.89 105.99 48.03 110.89 ;
      RECT  47.18 105.08 47.61 105.51 ;
      RECT  46.77 105.99 46.91 110.87 ;
      RECT  47.89 105.64 48.24 105.99 ;
      RECT  46.56 105.64 46.91 105.99 ;
      RECT  46.77 104.99 46.91 105.64 ;
      RECT  47.89 104.99 48.03 105.64 ;
      RECT  47.18 110.2 47.61 110.63 ;
      RECT  47.89 114.85 48.03 109.95 ;
      RECT  47.18 115.76 47.61 115.33 ;
      RECT  46.77 114.85 46.91 109.97 ;
      RECT  47.89 115.2 48.24 114.85 ;
      RECT  46.56 115.2 46.91 114.85 ;
      RECT  46.77 115.85 46.91 115.2 ;
      RECT  47.89 115.85 48.03 115.2 ;
      RECT  47.18 110.64 47.61 110.21 ;
      RECT  47.89 116.25 48.03 121.15 ;
      RECT  47.18 115.34 47.61 115.77 ;
      RECT  46.77 116.25 46.91 121.13 ;
      RECT  47.89 115.9 48.24 116.25 ;
      RECT  46.56 115.9 46.91 116.25 ;
      RECT  46.77 115.25 46.91 115.9 ;
      RECT  47.89 115.25 48.03 115.9 ;
      RECT  47.18 120.46 47.61 120.89 ;
      RECT  46.77 23.21 46.91 120.68 ;
      RECT  47.89 23.21 48.03 120.68 ;
      RECT  50.49 32.77 50.63 27.87 ;
      RECT  49.78 33.68 50.21 33.25 ;
      RECT  49.37 32.77 49.51 27.89 ;
      RECT  50.49 33.12 50.84 32.77 ;
      RECT  49.16 33.12 49.51 32.77 ;
      RECT  49.37 33.77 49.51 33.12 ;
      RECT  50.49 33.77 50.63 33.12 ;
      RECT  49.78 28.56 50.21 28.13 ;
      RECT  53.09 32.77 53.23 27.87 ;
      RECT  52.38 33.68 52.81 33.25 ;
      RECT  51.97 32.77 52.11 27.89 ;
      RECT  53.09 33.12 53.44 32.77 ;
      RECT  51.76 33.12 52.11 32.77 ;
      RECT  51.97 33.77 52.11 33.12 ;
      RECT  53.09 33.77 53.23 33.12 ;
      RECT  52.38 28.56 52.81 28.13 ;
      RECT  49.37 33.47 49.51 28.34 ;
      RECT  50.49 33.47 50.63 28.34 ;
      RECT  51.97 33.47 52.11 28.34 ;
      RECT  53.09 33.47 53.23 28.34 ;
      RECT  50.49 23.91 50.63 28.81 ;
      RECT  49.78 23.0 50.21 23.43 ;
      RECT  49.37 23.91 49.51 28.79 ;
      RECT  50.49 23.56 50.84 23.91 ;
      RECT  49.16 23.56 49.51 23.91 ;
      RECT  49.37 22.91 49.51 23.56 ;
      RECT  50.49 22.91 50.63 23.56 ;
      RECT  49.78 28.12 50.21 28.55 ;
      RECT  53.09 23.91 53.23 28.81 ;
      RECT  52.38 23.0 52.81 23.43 ;
      RECT  51.97 23.91 52.11 28.79 ;
      RECT  53.09 23.56 53.44 23.91 ;
      RECT  51.76 23.56 52.11 23.91 ;
      RECT  51.97 22.91 52.11 23.56 ;
      RECT  53.09 22.91 53.23 23.56 ;
      RECT  52.38 28.12 52.81 28.55 ;
      RECT  49.37 23.21 49.51 28.34 ;
      RECT  50.49 23.21 50.63 28.34 ;
      RECT  51.97 23.21 52.11 28.34 ;
      RECT  53.09 23.21 53.23 28.34 ;
      RECT  50.49 116.25 50.63 121.15 ;
      RECT  49.78 115.34 50.21 115.77 ;
      RECT  49.37 116.25 49.51 121.13 ;
      RECT  50.49 115.9 50.84 116.25 ;
      RECT  49.16 115.9 49.51 116.25 ;
      RECT  49.37 115.25 49.51 115.9 ;
      RECT  50.49 115.25 50.63 115.9 ;
      RECT  49.78 120.46 50.21 120.89 ;
      RECT  53.09 116.25 53.23 121.15 ;
      RECT  52.38 115.34 52.81 115.77 ;
      RECT  51.97 116.25 52.11 121.13 ;
      RECT  53.09 115.9 53.44 116.25 ;
      RECT  51.76 115.9 52.11 116.25 ;
      RECT  51.97 115.25 52.11 115.9 ;
      RECT  53.09 115.25 53.23 115.9 ;
      RECT  52.38 120.46 52.81 120.89 ;
      RECT  49.37 115.55 49.51 120.68 ;
      RECT  50.49 115.55 50.63 120.68 ;
      RECT  51.97 115.55 52.11 120.68 ;
      RECT  53.09 115.55 53.23 120.68 ;
      RECT  45.29 23.91 45.43 28.81 ;
      RECT  44.58 23.0 45.01 23.43 ;
      RECT  44.17 23.91 44.31 28.79 ;
      RECT  45.29 23.56 45.64 23.91 ;
      RECT  43.96 23.56 44.31 23.91 ;
      RECT  44.17 22.91 44.31 23.56 ;
      RECT  45.29 22.91 45.43 23.56 ;
      RECT  44.58 28.12 45.01 28.55 ;
      RECT  45.29 32.77 45.43 27.87 ;
      RECT  44.58 33.68 45.01 33.25 ;
      RECT  44.17 32.77 44.31 27.89 ;
      RECT  45.29 33.12 45.64 32.77 ;
      RECT  43.96 33.12 44.31 32.77 ;
      RECT  44.17 33.77 44.31 33.12 ;
      RECT  45.29 33.77 45.43 33.12 ;
      RECT  44.58 28.56 45.01 28.13 ;
      RECT  45.29 34.17 45.43 39.07 ;
      RECT  44.58 33.26 45.01 33.69 ;
      RECT  44.17 34.17 44.31 39.05 ;
      RECT  45.29 33.82 45.64 34.17 ;
      RECT  43.96 33.82 44.31 34.17 ;
      RECT  44.17 33.17 44.31 33.82 ;
      RECT  45.29 33.17 45.43 33.82 ;
      RECT  44.58 38.38 45.01 38.81 ;
      RECT  45.29 43.03 45.43 38.13 ;
      RECT  44.58 43.94 45.01 43.51 ;
      RECT  44.17 43.03 44.31 38.15 ;
      RECT  45.29 43.38 45.64 43.03 ;
      RECT  43.96 43.38 44.31 43.03 ;
      RECT  44.17 44.03 44.31 43.38 ;
      RECT  45.29 44.03 45.43 43.38 ;
      RECT  44.58 38.82 45.01 38.39 ;
      RECT  45.29 44.43 45.43 49.33 ;
      RECT  44.58 43.52 45.01 43.95 ;
      RECT  44.17 44.43 44.31 49.31 ;
      RECT  45.29 44.08 45.64 44.43 ;
      RECT  43.96 44.08 44.31 44.43 ;
      RECT  44.17 43.43 44.31 44.08 ;
      RECT  45.29 43.43 45.43 44.08 ;
      RECT  44.58 48.64 45.01 49.07 ;
      RECT  45.29 53.29 45.43 48.39 ;
      RECT  44.58 54.2 45.01 53.77 ;
      RECT  44.17 53.29 44.31 48.41 ;
      RECT  45.29 53.64 45.64 53.29 ;
      RECT  43.96 53.64 44.31 53.29 ;
      RECT  44.17 54.29 44.31 53.64 ;
      RECT  45.29 54.29 45.43 53.64 ;
      RECT  44.58 49.08 45.01 48.65 ;
      RECT  45.29 54.69 45.43 59.59 ;
      RECT  44.58 53.78 45.01 54.21 ;
      RECT  44.17 54.69 44.31 59.57 ;
      RECT  45.29 54.34 45.64 54.69 ;
      RECT  43.96 54.34 44.31 54.69 ;
      RECT  44.17 53.69 44.31 54.34 ;
      RECT  45.29 53.69 45.43 54.34 ;
      RECT  44.58 58.9 45.01 59.33 ;
      RECT  45.29 63.55 45.43 58.65 ;
      RECT  44.58 64.46 45.01 64.03 ;
      RECT  44.17 63.55 44.31 58.67 ;
      RECT  45.29 63.9 45.64 63.55 ;
      RECT  43.96 63.9 44.31 63.55 ;
      RECT  44.17 64.55 44.31 63.9 ;
      RECT  45.29 64.55 45.43 63.9 ;
      RECT  44.58 59.34 45.01 58.91 ;
      RECT  45.29 64.95 45.43 69.85 ;
      RECT  44.58 64.04 45.01 64.47 ;
      RECT  44.17 64.95 44.31 69.83 ;
      RECT  45.29 64.6 45.64 64.95 ;
      RECT  43.96 64.6 44.31 64.95 ;
      RECT  44.17 63.95 44.31 64.6 ;
      RECT  45.29 63.95 45.43 64.6 ;
      RECT  44.58 69.16 45.01 69.59 ;
      RECT  45.29 73.81 45.43 68.91 ;
      RECT  44.58 74.72 45.01 74.29 ;
      RECT  44.17 73.81 44.31 68.93 ;
      RECT  45.29 74.16 45.64 73.81 ;
      RECT  43.96 74.16 44.31 73.81 ;
      RECT  44.17 74.81 44.31 74.16 ;
      RECT  45.29 74.81 45.43 74.16 ;
      RECT  44.58 69.6 45.01 69.17 ;
      RECT  45.29 75.21 45.43 80.11 ;
      RECT  44.58 74.3 45.01 74.73 ;
      RECT  44.17 75.21 44.31 80.09 ;
      RECT  45.29 74.86 45.64 75.21 ;
      RECT  43.96 74.86 44.31 75.21 ;
      RECT  44.17 74.21 44.31 74.86 ;
      RECT  45.29 74.21 45.43 74.86 ;
      RECT  44.58 79.42 45.01 79.85 ;
      RECT  45.29 84.07 45.43 79.17 ;
      RECT  44.58 84.98 45.01 84.55 ;
      RECT  44.17 84.07 44.31 79.19 ;
      RECT  45.29 84.42 45.64 84.07 ;
      RECT  43.96 84.42 44.31 84.07 ;
      RECT  44.17 85.07 44.31 84.42 ;
      RECT  45.29 85.07 45.43 84.42 ;
      RECT  44.58 79.86 45.01 79.43 ;
      RECT  45.29 85.47 45.43 90.37 ;
      RECT  44.58 84.56 45.01 84.99 ;
      RECT  44.17 85.47 44.31 90.35 ;
      RECT  45.29 85.12 45.64 85.47 ;
      RECT  43.96 85.12 44.31 85.47 ;
      RECT  44.17 84.47 44.31 85.12 ;
      RECT  45.29 84.47 45.43 85.12 ;
      RECT  44.58 89.68 45.01 90.11 ;
      RECT  45.29 94.33 45.43 89.43 ;
      RECT  44.58 95.24 45.01 94.81 ;
      RECT  44.17 94.33 44.31 89.45 ;
      RECT  45.29 94.68 45.64 94.33 ;
      RECT  43.96 94.68 44.31 94.33 ;
      RECT  44.17 95.33 44.31 94.68 ;
      RECT  45.29 95.33 45.43 94.68 ;
      RECT  44.58 90.12 45.01 89.69 ;
      RECT  45.29 95.73 45.43 100.63 ;
      RECT  44.58 94.82 45.01 95.25 ;
      RECT  44.17 95.73 44.31 100.61 ;
      RECT  45.29 95.38 45.64 95.73 ;
      RECT  43.96 95.38 44.31 95.73 ;
      RECT  44.17 94.73 44.31 95.38 ;
      RECT  45.29 94.73 45.43 95.38 ;
      RECT  44.58 99.94 45.01 100.37 ;
      RECT  45.29 104.59 45.43 99.69 ;
      RECT  44.58 105.5 45.01 105.07 ;
      RECT  44.17 104.59 44.31 99.71 ;
      RECT  45.29 104.94 45.64 104.59 ;
      RECT  43.96 104.94 44.31 104.59 ;
      RECT  44.17 105.59 44.31 104.94 ;
      RECT  45.29 105.59 45.43 104.94 ;
      RECT  44.58 100.38 45.01 99.95 ;
      RECT  45.29 105.99 45.43 110.89 ;
      RECT  44.58 105.08 45.01 105.51 ;
      RECT  44.17 105.99 44.31 110.87 ;
      RECT  45.29 105.64 45.64 105.99 ;
      RECT  43.96 105.64 44.31 105.99 ;
      RECT  44.17 104.99 44.31 105.64 ;
      RECT  45.29 104.99 45.43 105.64 ;
      RECT  44.58 110.2 45.01 110.63 ;
      RECT  45.29 114.85 45.43 109.95 ;
      RECT  44.58 115.76 45.01 115.33 ;
      RECT  44.17 114.85 44.31 109.97 ;
      RECT  45.29 115.2 45.64 114.85 ;
      RECT  43.96 115.2 44.31 114.85 ;
      RECT  44.17 115.85 44.31 115.2 ;
      RECT  45.29 115.85 45.43 115.2 ;
      RECT  44.58 110.64 45.01 110.21 ;
      RECT  45.29 116.25 45.43 121.15 ;
      RECT  44.58 115.34 45.01 115.77 ;
      RECT  44.17 116.25 44.31 121.13 ;
      RECT  45.29 115.9 45.64 116.25 ;
      RECT  43.96 115.9 44.31 116.25 ;
      RECT  44.17 115.25 44.31 115.9 ;
      RECT  45.29 115.25 45.43 115.9 ;
      RECT  44.58 120.46 45.01 120.89 ;
      RECT  44.17 23.21 44.31 120.68 ;
      RECT  45.29 23.21 45.43 120.68 ;
      RECT  55.69 23.91 55.83 28.81 ;
      RECT  54.98 23.0 55.41 23.43 ;
      RECT  54.57 23.91 54.71 28.79 ;
      RECT  55.69 23.56 56.04 23.91 ;
      RECT  54.36 23.56 54.71 23.91 ;
      RECT  54.57 22.91 54.71 23.56 ;
      RECT  55.69 22.91 55.83 23.56 ;
      RECT  54.98 28.12 55.41 28.55 ;
      RECT  55.69 32.77 55.83 27.87 ;
      RECT  54.98 33.68 55.41 33.25 ;
      RECT  54.57 32.77 54.71 27.89 ;
      RECT  55.69 33.12 56.04 32.77 ;
      RECT  54.36 33.12 54.71 32.77 ;
      RECT  54.57 33.77 54.71 33.12 ;
      RECT  55.69 33.77 55.83 33.12 ;
      RECT  54.98 28.56 55.41 28.13 ;
      RECT  55.69 34.17 55.83 39.07 ;
      RECT  54.98 33.26 55.41 33.69 ;
      RECT  54.57 34.17 54.71 39.05 ;
      RECT  55.69 33.82 56.04 34.17 ;
      RECT  54.36 33.82 54.71 34.17 ;
      RECT  54.57 33.17 54.71 33.82 ;
      RECT  55.69 33.17 55.83 33.82 ;
      RECT  54.98 38.38 55.41 38.81 ;
      RECT  55.69 43.03 55.83 38.13 ;
      RECT  54.98 43.94 55.41 43.51 ;
      RECT  54.57 43.03 54.71 38.15 ;
      RECT  55.69 43.38 56.04 43.03 ;
      RECT  54.36 43.38 54.71 43.03 ;
      RECT  54.57 44.03 54.71 43.38 ;
      RECT  55.69 44.03 55.83 43.38 ;
      RECT  54.98 38.82 55.41 38.39 ;
      RECT  55.69 44.43 55.83 49.33 ;
      RECT  54.98 43.52 55.41 43.95 ;
      RECT  54.57 44.43 54.71 49.31 ;
      RECT  55.69 44.08 56.04 44.43 ;
      RECT  54.36 44.08 54.71 44.43 ;
      RECT  54.57 43.43 54.71 44.08 ;
      RECT  55.69 43.43 55.83 44.08 ;
      RECT  54.98 48.64 55.41 49.07 ;
      RECT  55.69 53.29 55.83 48.39 ;
      RECT  54.98 54.2 55.41 53.77 ;
      RECT  54.57 53.29 54.71 48.41 ;
      RECT  55.69 53.64 56.04 53.29 ;
      RECT  54.36 53.64 54.71 53.29 ;
      RECT  54.57 54.29 54.71 53.64 ;
      RECT  55.69 54.29 55.83 53.64 ;
      RECT  54.98 49.08 55.41 48.65 ;
      RECT  55.69 54.69 55.83 59.59 ;
      RECT  54.98 53.78 55.41 54.21 ;
      RECT  54.57 54.69 54.71 59.57 ;
      RECT  55.69 54.34 56.04 54.69 ;
      RECT  54.36 54.34 54.71 54.69 ;
      RECT  54.57 53.69 54.71 54.34 ;
      RECT  55.69 53.69 55.83 54.34 ;
      RECT  54.98 58.9 55.41 59.33 ;
      RECT  55.69 63.55 55.83 58.65 ;
      RECT  54.98 64.46 55.41 64.03 ;
      RECT  54.57 63.55 54.71 58.67 ;
      RECT  55.69 63.9 56.04 63.55 ;
      RECT  54.36 63.9 54.71 63.55 ;
      RECT  54.57 64.55 54.71 63.9 ;
      RECT  55.69 64.55 55.83 63.9 ;
      RECT  54.98 59.34 55.41 58.91 ;
      RECT  55.69 64.95 55.83 69.85 ;
      RECT  54.98 64.04 55.41 64.47 ;
      RECT  54.57 64.95 54.71 69.83 ;
      RECT  55.69 64.6 56.04 64.95 ;
      RECT  54.36 64.6 54.71 64.95 ;
      RECT  54.57 63.95 54.71 64.6 ;
      RECT  55.69 63.95 55.83 64.6 ;
      RECT  54.98 69.16 55.41 69.59 ;
      RECT  55.69 73.81 55.83 68.91 ;
      RECT  54.98 74.72 55.41 74.29 ;
      RECT  54.57 73.81 54.71 68.93 ;
      RECT  55.69 74.16 56.04 73.81 ;
      RECT  54.36 74.16 54.71 73.81 ;
      RECT  54.57 74.81 54.71 74.16 ;
      RECT  55.69 74.81 55.83 74.16 ;
      RECT  54.98 69.6 55.41 69.17 ;
      RECT  55.69 75.21 55.83 80.11 ;
      RECT  54.98 74.3 55.41 74.73 ;
      RECT  54.57 75.21 54.71 80.09 ;
      RECT  55.69 74.86 56.04 75.21 ;
      RECT  54.36 74.86 54.71 75.21 ;
      RECT  54.57 74.21 54.71 74.86 ;
      RECT  55.69 74.21 55.83 74.86 ;
      RECT  54.98 79.42 55.41 79.85 ;
      RECT  55.69 84.07 55.83 79.17 ;
      RECT  54.98 84.98 55.41 84.55 ;
      RECT  54.57 84.07 54.71 79.19 ;
      RECT  55.69 84.42 56.04 84.07 ;
      RECT  54.36 84.42 54.71 84.07 ;
      RECT  54.57 85.07 54.71 84.42 ;
      RECT  55.69 85.07 55.83 84.42 ;
      RECT  54.98 79.86 55.41 79.43 ;
      RECT  55.69 85.47 55.83 90.37 ;
      RECT  54.98 84.56 55.41 84.99 ;
      RECT  54.57 85.47 54.71 90.35 ;
      RECT  55.69 85.12 56.04 85.47 ;
      RECT  54.36 85.12 54.71 85.47 ;
      RECT  54.57 84.47 54.71 85.12 ;
      RECT  55.69 84.47 55.83 85.12 ;
      RECT  54.98 89.68 55.41 90.11 ;
      RECT  55.69 94.33 55.83 89.43 ;
      RECT  54.98 95.24 55.41 94.81 ;
      RECT  54.57 94.33 54.71 89.45 ;
      RECT  55.69 94.68 56.04 94.33 ;
      RECT  54.36 94.68 54.71 94.33 ;
      RECT  54.57 95.33 54.71 94.68 ;
      RECT  55.69 95.33 55.83 94.68 ;
      RECT  54.98 90.12 55.41 89.69 ;
      RECT  55.69 95.73 55.83 100.63 ;
      RECT  54.98 94.82 55.41 95.25 ;
      RECT  54.57 95.73 54.71 100.61 ;
      RECT  55.69 95.38 56.04 95.73 ;
      RECT  54.36 95.38 54.71 95.73 ;
      RECT  54.57 94.73 54.71 95.38 ;
      RECT  55.69 94.73 55.83 95.38 ;
      RECT  54.98 99.94 55.41 100.37 ;
      RECT  55.69 104.59 55.83 99.69 ;
      RECT  54.98 105.5 55.41 105.07 ;
      RECT  54.57 104.59 54.71 99.71 ;
      RECT  55.69 104.94 56.04 104.59 ;
      RECT  54.36 104.94 54.71 104.59 ;
      RECT  54.57 105.59 54.71 104.94 ;
      RECT  55.69 105.59 55.83 104.94 ;
      RECT  54.98 100.38 55.41 99.95 ;
      RECT  55.69 105.99 55.83 110.89 ;
      RECT  54.98 105.08 55.41 105.51 ;
      RECT  54.57 105.99 54.71 110.87 ;
      RECT  55.69 105.64 56.04 105.99 ;
      RECT  54.36 105.64 54.71 105.99 ;
      RECT  54.57 104.99 54.71 105.64 ;
      RECT  55.69 104.99 55.83 105.64 ;
      RECT  54.98 110.2 55.41 110.63 ;
      RECT  55.69 114.85 55.83 109.95 ;
      RECT  54.98 115.76 55.41 115.33 ;
      RECT  54.57 114.85 54.71 109.97 ;
      RECT  55.69 115.2 56.04 114.85 ;
      RECT  54.36 115.2 54.71 114.85 ;
      RECT  54.57 115.85 54.71 115.2 ;
      RECT  55.69 115.85 55.83 115.2 ;
      RECT  54.98 110.64 55.41 110.21 ;
      RECT  55.69 116.25 55.83 121.15 ;
      RECT  54.98 115.34 55.41 115.77 ;
      RECT  54.57 116.25 54.71 121.13 ;
      RECT  55.69 115.9 56.04 116.25 ;
      RECT  54.36 115.9 54.71 116.25 ;
      RECT  54.57 115.25 54.71 115.9 ;
      RECT  55.69 115.25 55.83 115.9 ;
      RECT  54.98 120.46 55.41 120.89 ;
      RECT  54.57 23.21 54.71 120.68 ;
      RECT  55.69 23.21 55.83 120.68 ;
      RECT  46.77 23.21 46.91 120.68 ;
      RECT  47.89 23.21 48.03 120.68 ;
      RECT  49.37 23.21 49.51 120.68 ;
      RECT  50.49 23.21 50.63 120.68 ;
      RECT  51.97 23.21 52.11 120.68 ;
      RECT  53.09 23.21 53.23 120.68 ;
      RECT  46.64 14.23 46.78 21.23 ;
      RECT  47.92 14.23 48.06 21.23 ;
      RECT  49.24 14.23 49.38 21.23 ;
      RECT  50.52 14.23 50.66 21.23 ;
      RECT  51.84 14.23 51.98 21.23 ;
      RECT  53.12 14.23 53.26 21.23 ;
      RECT  46.64 14.23 46.78 21.23 ;
      RECT  47.92 14.23 48.06 21.23 ;
      RECT  49.24 14.23 49.38 21.23 ;
      RECT  50.52 14.23 50.66 21.23 ;
      RECT  51.84 14.23 51.98 21.23 ;
      RECT  53.12 14.23 53.26 21.23 ;
      RECT  51.26 9.47 51.4 12.7 ;
      RECT  50.15 7.59 50.29 9.76 ;
      RECT  51.26 9.14 51.72 9.47 ;
      RECT  51.26 7.59 51.4 9.14 ;
      RECT  51.95 7.57 52.4 8.02 ;
      RECT  50.15 10.09 50.29 12.7 ;
      RECT  50.15 9.76 50.48 10.09 ;
      RECT  51.81 12.03 52.26 12.48 ;
      RECT  53.86 9.47 54.0 12.7 ;
      RECT  52.75 7.59 52.89 9.76 ;
      RECT  53.86 9.14 54.32 9.47 ;
      RECT  53.86 7.59 54.0 9.14 ;
      RECT  54.55 7.57 55.0 8.02 ;
      RECT  52.75 10.09 52.89 12.7 ;
      RECT  52.75 9.76 53.08 10.09 ;
      RECT  54.41 12.03 54.86 12.48 ;
      RECT  50.15 9.76 50.48 10.09 ;
      RECT  51.26 9.14 51.72 9.47 ;
      RECT  52.75 9.76 53.08 10.09 ;
      RECT  53.86 9.14 54.32 9.47 ;
      RECT  46.64 21.23 46.78 14.23 ;
      RECT  47.92 21.23 48.06 14.23 ;
      RECT  49.24 21.23 49.38 14.23 ;
      RECT  50.52 21.23 50.66 14.23 ;
      RECT  51.84 21.23 51.98 14.23 ;
      RECT  53.12 21.23 53.26 14.23 ;
      RECT  3.44 35.7 3.9 36.16 ;
      RECT  4.1 41.04 4.56 41.5 ;
      RECT  3.44 66.48 3.9 66.94 ;
      RECT  4.1 71.82 4.56 72.28 ;
      RECT  0.16 33.47 0.3 84.77 ;
      RECT  0.82 33.47 0.96 84.77 ;
      RECT  1.48 33.47 1.62 84.77 ;
      RECT  2.14 33.47 2.28 84.77 ;
      RECT  34.585 33.47 34.725 115.55 ;
      RECT  0.16 33.47 0.3 84.77 ;
      RECT  0.82 33.47 0.96 84.77 ;
      RECT  1.48 33.47 1.62 84.77 ;
      RECT  2.14 33.47 2.28 84.77 ;
      RECT  34.09 31.885 34.23 32.025 ;
      RECT  0.16 33.47 0.3 84.77 ;
      RECT  0.82 33.47 0.96 84.77 ;
      RECT  1.48 33.47 1.62 84.77 ;
      RECT  2.14 33.47 2.28 84.77 ;
      RECT  37.63 0.0 37.77 23.21 ;
      RECT  39.27 0.0 39.41 23.21 ;
      RECT  38.45 0.0 38.59 23.21 ;
      RECT  40.09 0.0 40.23 23.21 ;
      RECT  -54.22 -8.38 -53.88 -8.06 ;
      RECT  -55.0 -9.2 -54.69 -8.88 ;
      RECT  -45.32 -8.69 -45.0 -8.37 ;
      RECT  -54.22 -8.38 -53.88 -8.06 ;
      RECT  -32.755 -10.195 -32.615 -10.055 ;
      RECT  -36.52 -7.52 -36.38 -7.38 ;
      RECT  -55.0 -9.2 -54.69 -8.88 ;
      RECT  -54.22 -4.86 -53.88 -5.18 ;
      RECT  -55.0 -4.04 -54.69 -4.36 ;
      RECT  -45.32 -4.55 -45.0 -4.87 ;
      RECT  -54.22 -4.86 -53.88 -5.18 ;
      RECT  -32.755 -3.045 -32.615 -3.185 ;
      RECT  -36.52 -5.72 -36.38 -5.86 ;
      RECT  -55.0 -4.04 -54.69 -4.36 ;
      RECT  -54.22 -8.38 -53.88 -8.06 ;
      RECT  -54.22 -5.18 -53.88 -4.86 ;
      RECT  -32.755 -10.195 -32.615 -10.055 ;
      RECT  -36.52 -7.52 -36.38 -7.38 ;
      RECT  -32.755 -3.185 -32.615 -3.045 ;
      RECT  -36.52 -5.86 -36.38 -5.72 ;
      RECT  -55.0 -10.71 -54.86 -2.53 ;
      RECT  -40.955 23.21 -41.095 27.305 ;
      RECT  -54.03 23.21 -54.17 94.505 ;
      RECT  -54.22 -8.38 -53.88 -8.06 ;
      RECT  -54.22 -5.18 -53.88 -4.86 ;
      RECT  -24.34 -8.84 -24.2 -8.7 ;
      RECT  -41.095 23.21 -40.955 27.305 ;
      RECT  -18.795 20.0 -1.32 20.14 ;
      RECT  -16.505 7.475 -1.32 7.615 ;
      RECT  -16.66 11.82 -1.32 11.96 ;
      RECT  -11.815 3.665 -1.32 3.805 ;
      RECT  -7.135 -8.895 -1.32 -8.755 ;
      RECT  -12.8 102.34 -12.46 102.66 ;
      RECT  -13.58 101.52 -13.27 101.84 ;
      RECT  -3.9 102.03 -3.58 102.35 ;
      RECT  -12.8 105.86 -12.46 105.54 ;
      RECT  -13.58 106.68 -13.27 106.36 ;
      RECT  -3.9 106.17 -3.58 105.85 ;
      RECT  -12.8 110.52 -12.46 110.84 ;
      RECT  -13.58 109.7 -13.27 110.02 ;
      RECT  -3.9 110.21 -3.58 110.53 ;
      RECT  -12.8 114.04 -12.46 113.72 ;
      RECT  -13.58 114.86 -13.27 114.54 ;
      RECT  -3.9 114.35 -3.58 114.03 ;
      RECT  -12.8 102.34 -12.46 102.66 ;
      RECT  -12.8 105.54 -12.46 105.86 ;
      RECT  -12.8 110.52 -12.46 110.84 ;
      RECT  -12.8 113.72 -12.46 114.04 ;
      RECT  -3.9 102.03 -3.58 102.35 ;
      RECT  -3.9 105.85 -3.58 106.17 ;
      RECT  -3.9 110.21 -3.58 110.53 ;
      RECT  -3.9 114.03 -3.58 114.35 ;
      RECT  12.62 -8.38 12.96 -8.06 ;
      RECT  11.84 -9.2 12.15 -8.88 ;
      RECT  21.52 -8.69 21.84 -8.37 ;
      RECT  25.33 -8.38 25.67 -8.06 ;
      RECT  24.55 -9.2 24.86 -8.88 ;
      RECT  34.23 -8.69 34.55 -8.37 ;
      RECT  12.62 -8.38 12.96 -8.06 ;
      RECT  25.33 -8.38 25.67 -8.06 ;
      RECT  21.52 -8.69 21.84 -8.37 ;
      RECT  34.23 -8.69 34.55 -8.37 ;
   LAYER  m3 ;
      RECT  49.7 33.17 50.3 33.77 ;
      RECT  49.7 38.29 50.3 38.89 ;
      RECT  49.7 44.03 50.3 43.43 ;
      RECT  49.7 38.91 50.3 38.31 ;
      RECT  49.7 43.43 50.3 44.03 ;
      RECT  49.7 48.55 50.3 49.15 ;
      RECT  49.7 54.29 50.3 53.69 ;
      RECT  49.7 49.17 50.3 48.57 ;
      RECT  49.7 53.69 50.3 54.29 ;
      RECT  49.7 58.81 50.3 59.41 ;
      RECT  49.7 64.55 50.3 63.95 ;
      RECT  49.7 59.43 50.3 58.83 ;
      RECT  49.7 63.95 50.3 64.55 ;
      RECT  49.7 69.07 50.3 69.67 ;
      RECT  49.7 74.81 50.3 74.21 ;
      RECT  49.7 69.69 50.3 69.09 ;
      RECT  49.7 74.21 50.3 74.81 ;
      RECT  49.7 79.33 50.3 79.93 ;
      RECT  49.7 85.07 50.3 84.47 ;
      RECT  49.7 79.95 50.3 79.35 ;
      RECT  49.7 84.47 50.3 85.07 ;
      RECT  49.7 89.59 50.3 90.19 ;
      RECT  49.7 95.33 50.3 94.73 ;
      RECT  49.7 90.21 50.3 89.61 ;
      RECT  49.7 94.73 50.3 95.33 ;
      RECT  49.7 99.85 50.3 100.45 ;
      RECT  49.7 105.59 50.3 104.99 ;
      RECT  49.7 100.47 50.3 99.87 ;
      RECT  49.7 104.99 50.3 105.59 ;
      RECT  49.7 110.11 50.3 110.71 ;
      RECT  49.7 115.85 50.3 115.25 ;
      RECT  49.7 110.73 50.3 110.13 ;
      RECT  52.3 33.17 52.9 33.77 ;
      RECT  52.3 38.29 52.9 38.89 ;
      RECT  52.3 44.03 52.9 43.43 ;
      RECT  52.3 38.91 52.9 38.31 ;
      RECT  52.3 43.43 52.9 44.03 ;
      RECT  52.3 48.55 52.9 49.15 ;
      RECT  52.3 54.29 52.9 53.69 ;
      RECT  52.3 49.17 52.9 48.57 ;
      RECT  52.3 53.69 52.9 54.29 ;
      RECT  52.3 58.81 52.9 59.41 ;
      RECT  52.3 64.55 52.9 63.95 ;
      RECT  52.3 59.43 52.9 58.83 ;
      RECT  52.3 63.95 52.9 64.55 ;
      RECT  52.3 69.07 52.9 69.67 ;
      RECT  52.3 74.81 52.9 74.21 ;
      RECT  52.3 69.69 52.9 69.09 ;
      RECT  52.3 74.21 52.9 74.81 ;
      RECT  52.3 79.33 52.9 79.93 ;
      RECT  52.3 85.07 52.9 84.47 ;
      RECT  52.3 79.95 52.9 79.35 ;
      RECT  52.3 84.47 52.9 85.07 ;
      RECT  52.3 89.59 52.9 90.19 ;
      RECT  52.3 95.33 52.9 94.73 ;
      RECT  52.3 90.21 52.9 89.61 ;
      RECT  52.3 94.73 52.9 95.33 ;
      RECT  52.3 99.85 52.9 100.45 ;
      RECT  52.3 105.59 52.9 104.99 ;
      RECT  52.3 100.47 52.9 99.87 ;
      RECT  52.3 104.99 52.9 105.59 ;
      RECT  52.3 110.11 52.9 110.71 ;
      RECT  52.3 115.85 52.9 115.25 ;
      RECT  52.3 110.73 52.9 110.13 ;
      RECT  47.1 22.91 47.7 23.51 ;
      RECT  47.1 28.03 47.7 28.63 ;
      RECT  47.1 33.77 47.7 33.17 ;
      RECT  47.1 28.65 47.7 28.05 ;
      RECT  47.1 33.17 47.7 33.77 ;
      RECT  47.1 38.29 47.7 38.89 ;
      RECT  47.1 44.03 47.7 43.43 ;
      RECT  47.1 38.91 47.7 38.31 ;
      RECT  47.1 43.43 47.7 44.03 ;
      RECT  47.1 48.55 47.7 49.15 ;
      RECT  47.1 54.29 47.7 53.69 ;
      RECT  47.1 49.17 47.7 48.57 ;
      RECT  47.1 53.69 47.7 54.29 ;
      RECT  47.1 58.81 47.7 59.41 ;
      RECT  47.1 64.55 47.7 63.95 ;
      RECT  47.1 59.43 47.7 58.83 ;
      RECT  47.1 63.95 47.7 64.55 ;
      RECT  47.1 69.07 47.7 69.67 ;
      RECT  47.1 74.81 47.7 74.21 ;
      RECT  47.1 69.69 47.7 69.09 ;
      RECT  47.1 74.21 47.7 74.81 ;
      RECT  47.1 79.33 47.7 79.93 ;
      RECT  47.1 85.07 47.7 84.47 ;
      RECT  47.1 79.95 47.7 79.35 ;
      RECT  47.1 84.47 47.7 85.07 ;
      RECT  47.1 89.59 47.7 90.19 ;
      RECT  47.1 95.33 47.7 94.73 ;
      RECT  47.1 90.21 47.7 89.61 ;
      RECT  47.1 94.73 47.7 95.33 ;
      RECT  47.1 99.85 47.7 100.45 ;
      RECT  47.1 105.59 47.7 104.99 ;
      RECT  47.1 100.47 47.7 99.87 ;
      RECT  47.1 104.99 47.7 105.59 ;
      RECT  47.1 110.11 47.7 110.71 ;
      RECT  47.1 115.85 47.7 115.25 ;
      RECT  47.1 110.73 47.7 110.13 ;
      RECT  47.1 115.25 47.7 115.85 ;
      RECT  47.1 120.37 47.7 120.97 ;
      RECT  47.09 28.075 47.61 28.595 ;
      RECT  47.09 120.415 47.61 120.935 ;
      RECT  47.09 22.955 47.61 23.475 ;
      RECT  47.09 115.295 47.61 115.815 ;
      RECT  49.7 33.77 50.3 33.17 ;
      RECT  49.7 28.65 50.3 28.05 ;
      RECT  52.3 33.77 52.9 33.17 ;
      RECT  52.3 28.65 52.9 28.05 ;
      RECT  49.7 22.91 50.3 23.51 ;
      RECT  49.7 28.03 50.3 28.63 ;
      RECT  52.3 22.91 52.9 23.51 ;
      RECT  52.3 28.03 52.9 28.63 ;
      RECT  49.7 115.25 50.3 115.85 ;
      RECT  49.7 120.37 50.3 120.97 ;
      RECT  52.3 115.25 52.9 115.85 ;
      RECT  52.3 120.37 52.9 120.97 ;
      RECT  44.5 22.91 45.1 23.51 ;
      RECT  44.5 28.03 45.1 28.63 ;
      RECT  44.5 33.77 45.1 33.17 ;
      RECT  44.5 28.65 45.1 28.05 ;
      RECT  44.5 33.17 45.1 33.77 ;
      RECT  44.5 38.29 45.1 38.89 ;
      RECT  44.5 44.03 45.1 43.43 ;
      RECT  44.5 38.91 45.1 38.31 ;
      RECT  44.5 43.43 45.1 44.03 ;
      RECT  44.5 48.55 45.1 49.15 ;
      RECT  44.5 54.29 45.1 53.69 ;
      RECT  44.5 49.17 45.1 48.57 ;
      RECT  44.5 53.69 45.1 54.29 ;
      RECT  44.5 58.81 45.1 59.41 ;
      RECT  44.5 64.55 45.1 63.95 ;
      RECT  44.5 59.43 45.1 58.83 ;
      RECT  44.5 63.95 45.1 64.55 ;
      RECT  44.5 69.07 45.1 69.67 ;
      RECT  44.5 74.81 45.1 74.21 ;
      RECT  44.5 69.69 45.1 69.09 ;
      RECT  44.5 74.21 45.1 74.81 ;
      RECT  44.5 79.33 45.1 79.93 ;
      RECT  44.5 85.07 45.1 84.47 ;
      RECT  44.5 79.95 45.1 79.35 ;
      RECT  44.5 84.47 45.1 85.07 ;
      RECT  44.5 89.59 45.1 90.19 ;
      RECT  44.5 95.33 45.1 94.73 ;
      RECT  44.5 90.21 45.1 89.61 ;
      RECT  44.5 94.73 45.1 95.33 ;
      RECT  44.5 99.85 45.1 100.45 ;
      RECT  44.5 105.59 45.1 104.99 ;
      RECT  44.5 100.47 45.1 99.87 ;
      RECT  44.5 104.99 45.1 105.59 ;
      RECT  44.5 110.11 45.1 110.71 ;
      RECT  44.5 115.85 45.1 115.25 ;
      RECT  44.5 110.73 45.1 110.13 ;
      RECT  44.5 115.25 45.1 115.85 ;
      RECT  44.5 120.37 45.1 120.97 ;
      RECT  54.9 22.91 55.5 23.51 ;
      RECT  54.9 28.03 55.5 28.63 ;
      RECT  54.9 33.77 55.5 33.17 ;
      RECT  54.9 28.65 55.5 28.05 ;
      RECT  54.9 33.17 55.5 33.77 ;
      RECT  54.9 38.29 55.5 38.89 ;
      RECT  54.9 44.03 55.5 43.43 ;
      RECT  54.9 38.91 55.5 38.31 ;
      RECT  54.9 43.43 55.5 44.03 ;
      RECT  54.9 48.55 55.5 49.15 ;
      RECT  54.9 54.29 55.5 53.69 ;
      RECT  54.9 49.17 55.5 48.57 ;
      RECT  54.9 53.69 55.5 54.29 ;
      RECT  54.9 58.81 55.5 59.41 ;
      RECT  54.9 64.55 55.5 63.95 ;
      RECT  54.9 59.43 55.5 58.83 ;
      RECT  54.9 63.95 55.5 64.55 ;
      RECT  54.9 69.07 55.5 69.67 ;
      RECT  54.9 74.81 55.5 74.21 ;
      RECT  54.9 69.69 55.5 69.09 ;
      RECT  54.9 74.21 55.5 74.81 ;
      RECT  54.9 79.33 55.5 79.93 ;
      RECT  54.9 85.07 55.5 84.47 ;
      RECT  54.9 79.95 55.5 79.35 ;
      RECT  54.9 84.47 55.5 85.07 ;
      RECT  54.9 89.59 55.5 90.19 ;
      RECT  54.9 95.33 55.5 94.73 ;
      RECT  54.9 90.21 55.5 89.61 ;
      RECT  54.9 94.73 55.5 95.33 ;
      RECT  54.9 99.85 55.5 100.45 ;
      RECT  54.9 105.59 55.5 104.99 ;
      RECT  54.9 100.47 55.5 99.87 ;
      RECT  54.9 104.99 55.5 105.59 ;
      RECT  54.9 110.11 55.5 110.71 ;
      RECT  54.9 115.85 55.5 115.25 ;
      RECT  54.9 110.73 55.5 110.13 ;
      RECT  54.9 115.25 55.5 115.85 ;
      RECT  54.9 120.37 55.5 120.97 ;
      RECT  54.89 89.645 55.41 90.165 ;
      RECT  54.89 69.115 55.41 69.635 ;
      RECT  54.89 28.075 55.41 28.595 ;
      RECT  44.49 48.605 45.01 49.125 ;
      RECT  54.89 99.905 55.41 100.425 ;
      RECT  44.49 89.635 45.01 90.155 ;
      RECT  44.49 79.375 45.01 79.895 ;
      RECT  44.49 58.855 45.01 59.375 ;
      RECT  54.89 58.865 55.41 59.385 ;
      RECT  54.89 38.335 55.41 38.855 ;
      RECT  44.49 38.335 45.01 38.855 ;
      RECT  44.49 69.125 45.01 69.645 ;
      RECT  54.89 89.635 55.41 90.155 ;
      RECT  54.89 38.345 55.41 38.865 ;
      RECT  54.89 99.895 55.41 100.415 ;
      RECT  44.49 120.415 45.01 120.935 ;
      RECT  54.89 110.155 55.41 110.675 ;
      RECT  47.09 120.415 47.61 120.935 ;
      RECT  44.49 48.595 45.01 49.115 ;
      RECT  44.49 28.075 45.01 28.595 ;
      RECT  54.89 48.595 55.41 49.115 ;
      RECT  44.49 38.345 45.01 38.865 ;
      RECT  44.49 99.895 45.01 100.415 ;
      RECT  49.69 120.415 50.21 120.935 ;
      RECT  52.29 28.075 52.81 28.595 ;
      RECT  44.49 110.155 45.01 110.675 ;
      RECT  44.49 58.865 45.01 59.385 ;
      RECT  44.49 28.085 45.01 28.605 ;
      RECT  54.89 69.125 55.41 69.645 ;
      RECT  54.89 79.375 55.41 79.895 ;
      RECT  54.89 58.855 55.41 59.375 ;
      RECT  54.89 110.165 55.41 110.685 ;
      RECT  54.89 120.415 55.41 120.935 ;
      RECT  54.89 28.085 55.41 28.605 ;
      RECT  44.49 79.385 45.01 79.905 ;
      RECT  49.69 28.075 50.21 28.595 ;
      RECT  54.89 79.385 55.41 79.905 ;
      RECT  44.49 69.115 45.01 69.635 ;
      RECT  47.09 28.075 47.61 28.595 ;
      RECT  52.29 120.415 52.81 120.935 ;
      RECT  44.49 99.905 45.01 100.425 ;
      RECT  44.49 89.645 45.01 90.165 ;
      RECT  54.89 48.605 55.41 49.125 ;
      RECT  44.49 110.165 45.01 110.685 ;
      RECT  44.49 33.205 45.01 33.725 ;
      RECT  57.09 116.38 57.61 116.9 ;
      RECT  44.49 105.025 45.01 105.545 ;
      RECT  44.49 74.245 45.01 74.765 ;
      RECT  42.29 24.04 42.81 24.56 ;
      RECT  44.49 115.295 45.01 115.815 ;
      RECT  42.29 116.38 42.81 116.9 ;
      RECT  44.49 22.955 45.01 23.475 ;
      RECT  57.09 24.04 57.61 24.56 ;
      RECT  44.49 94.775 45.01 95.295 ;
      RECT  54.89 84.505 55.41 85.025 ;
      RECT  44.49 105.035 45.01 105.555 ;
      RECT  44.49 63.995 45.01 64.515 ;
      RECT  44.49 84.505 45.01 85.025 ;
      RECT  49.69 115.295 50.21 115.815 ;
      RECT  54.89 63.995 55.41 64.515 ;
      RECT  47.09 22.955 47.61 23.475 ;
      RECT  54.89 43.475 55.41 43.995 ;
      RECT  54.89 115.285 55.41 115.805 ;
      RECT  54.89 115.295 55.41 115.815 ;
      RECT  44.49 53.735 45.01 54.255 ;
      RECT  54.89 84.515 55.41 85.035 ;
      RECT  54.89 105.035 55.41 105.555 ;
      RECT  52.29 22.955 52.81 23.475 ;
      RECT  54.89 74.245 55.41 74.765 ;
      RECT  47.09 115.295 47.61 115.815 ;
      RECT  54.89 43.465 55.41 43.985 ;
      RECT  44.49 94.765 45.01 95.285 ;
      RECT  44.49 33.215 45.01 33.735 ;
      RECT  52.29 115.295 52.81 115.815 ;
      RECT  54.89 94.775 55.41 95.295 ;
      RECT  54.89 53.725 55.41 54.245 ;
      RECT  54.89 74.255 55.41 74.775 ;
      RECT  54.89 105.025 55.41 105.545 ;
      RECT  44.49 43.475 45.01 43.995 ;
      RECT  54.89 63.985 55.41 64.505 ;
      RECT  54.89 33.205 55.41 33.725 ;
      RECT  54.89 22.955 55.41 23.475 ;
      RECT  44.49 74.255 45.01 74.775 ;
      RECT  54.89 33.215 55.41 33.735 ;
      RECT  49.69 22.955 50.21 23.475 ;
      RECT  44.49 43.465 45.01 43.985 ;
      RECT  44.49 115.285 45.01 115.805 ;
      RECT  44.49 63.985 45.01 64.505 ;
      RECT  54.89 94.765 55.41 95.285 ;
      RECT  44.49 84.515 45.01 85.035 ;
      RECT  44.49 53.725 45.01 54.245 ;
      RECT  54.89 53.735 55.41 54.255 ;
      RECT  47.885 20.5 48.405 21.02 ;
      RECT  50.485 20.5 51.005 21.02 ;
      RECT  53.085 20.5 53.605 21.02 ;
      RECT  50.485 20.5 51.005 21.02 ;
      RECT  53.085 20.5 53.605 21.02 ;
      RECT  47.885 20.5 48.405 21.02 ;
      RECT  51.9 7.55 52.42 8.05 ;
      RECT  51.75 12.0 52.28 12.5 ;
      RECT  54.5 7.55 55.02 8.05 ;
      RECT  54.35 12.0 54.88 12.5 ;
      RECT  52.99 11.995 53.51 12.515 ;
      RECT  50.39 11.995 50.91 12.515 ;
      RECT  50.39 7.535 50.91 8.055 ;
      RECT  52.99 7.535 53.51 8.055 ;
      RECT  57.81 5.545 58.33 6.065 ;
      RECT  55.21 5.545 55.73 6.065 ;
      RECT  55.21 -0.265 55.73 0.255 ;
      RECT  57.81 -0.265 58.33 0.255 ;
      RECT  50.39 12.515 50.91 11.995 ;
      RECT  53.085 21.02 53.605 20.5 ;
      RECT  55.21 6.065 55.73 5.545 ;
      RECT  57.81 6.065 58.33 5.545 ;
      RECT  47.885 21.02 48.405 20.5 ;
      RECT  52.99 12.515 53.51 11.995 ;
      RECT  50.485 21.02 51.005 20.5 ;
      RECT  50.39 8.055 50.91 7.535 ;
      RECT  55.21 0.255 55.73 -0.265 ;
      RECT  52.99 8.055 53.51 7.535 ;
      RECT  57.81 0.255 58.33 -0.265 ;
      RECT  5.18 38.34 5.7 38.86 ;
      RECT  12.28 38.34 12.8 38.86 ;
      RECT  5.18 48.6 5.7 49.12 ;
      RECT  12.28 48.6 12.8 49.12 ;
      RECT  12.28 53.73 12.8 54.25 ;
      RECT  12.28 43.47 12.8 43.99 ;
      RECT  5.18 53.73 5.7 54.25 ;
      RECT  12.28 33.21 12.8 33.73 ;
      RECT  5.18 43.47 5.7 43.99 ;
      RECT  5.18 33.21 5.7 33.73 ;
      RECT  5.18 69.12 5.7 69.64 ;
      RECT  12.28 69.12 12.8 69.64 ;
      RECT  5.18 79.38 5.7 79.9 ;
      RECT  12.28 79.38 12.8 79.9 ;
      RECT  12.28 84.51 12.8 85.03 ;
      RECT  12.28 74.25 12.8 74.77 ;
      RECT  5.18 84.51 5.7 85.03 ;
      RECT  12.28 63.99 12.8 64.51 ;
      RECT  5.18 74.25 5.7 74.77 ;
      RECT  5.18 63.99 5.7 64.51 ;
      RECT  32.17 58.86 32.69 59.38 ;
      RECT  12.28 79.38 12.8 79.9 ;
      RECT  5.18 48.6 5.7 49.12 ;
      RECT  32.17 69.12 32.69 69.64 ;
      RECT  32.17 69.12 32.69 69.64 ;
      RECT  32.17 89.64 32.69 90.16 ;
      RECT  32.17 89.64 32.69 90.16 ;
      RECT  12.28 48.6 12.8 49.12 ;
      RECT  12.28 38.34 12.8 38.86 ;
      RECT  32.17 99.9 32.69 100.42 ;
      RECT  32.17 48.6 32.69 49.12 ;
      RECT  5.18 69.12 5.7 69.64 ;
      RECT  32.17 38.34 32.69 38.86 ;
      RECT  5.18 38.34 5.7 38.86 ;
      RECT  5.18 79.38 5.7 79.9 ;
      RECT  32.17 79.38 32.69 79.9 ;
      RECT  12.28 69.12 12.8 69.64 ;
      RECT  32.17 110.16 32.69 110.68 ;
      RECT  32.17 110.16 32.69 110.68 ;
      RECT  12.28 63.99 12.8 64.51 ;
      RECT  32.17 105.03 32.69 105.55 ;
      RECT  12.28 33.21 12.8 33.73 ;
      RECT  32.17 84.51 32.69 85.03 ;
      RECT  5.18 33.21 5.7 33.73 ;
      RECT  5.18 63.99 5.7 64.51 ;
      RECT  32.17 63.99 32.69 64.51 ;
      RECT  12.28 53.73 12.8 54.25 ;
      RECT  5.18 84.51 5.7 85.03 ;
      RECT  32.17 33.21 32.69 33.73 ;
      RECT  32.17 74.25 32.69 74.77 ;
      RECT  12.28 74.25 12.8 74.77 ;
      RECT  32.17 53.73 32.69 54.25 ;
      RECT  12.28 84.51 12.8 85.03 ;
      RECT  32.17 43.47 32.69 43.99 ;
      RECT  32.17 115.29 32.69 115.81 ;
      RECT  32.17 94.77 32.69 95.29 ;
      RECT  12.28 43.47 12.8 43.99 ;
      RECT  5.18 74.25 5.7 74.77 ;
      RECT  5.18 43.47 5.7 43.99 ;
      RECT  5.18 53.73 5.7 54.25 ;
      RECT  39.04 69.12 39.56 69.64 ;
      RECT  39.04 69.12 39.56 69.64 ;
      RECT  39.04 99.9 39.56 100.42 ;
      RECT  39.04 48.6 39.56 49.12 ;
      RECT  39.04 38.34 39.56 38.86 ;
      RECT  39.04 110.16 39.56 110.68 ;
      RECT  39.04 89.64 39.56 90.16 ;
      RECT  39.04 89.64 39.56 90.16 ;
      RECT  39.04 79.38 39.56 79.9 ;
      RECT  39.04 110.16 39.56 110.68 ;
      RECT  39.04 58.86 39.56 59.38 ;
      RECT  39.04 63.99 39.56 64.51 ;
      RECT  39.04 84.51 39.56 85.03 ;
      RECT  39.04 74.25 39.56 74.77 ;
      RECT  39.04 94.77 39.56 95.29 ;
      RECT  39.04 115.29 39.56 115.81 ;
      RECT  39.04 33.21 39.56 33.73 ;
      RECT  39.04 53.73 39.56 54.25 ;
      RECT  39.04 43.47 39.56 43.99 ;
      RECT  39.04 105.03 39.56 105.55 ;
      RECT  39.04 69.12 39.56 69.64 ;
      RECT  12.28 79.38 12.8 79.9 ;
      RECT  32.17 99.9 32.69 100.42 ;
      RECT  39.04 99.9 39.56 100.42 ;
      RECT  5.18 79.38 5.7 79.9 ;
      RECT  12.28 48.6 12.8 49.12 ;
      RECT  32.17 38.34 32.69 38.86 ;
      RECT  12.28 38.34 12.8 38.86 ;
      RECT  12.28 69.12 12.8 69.64 ;
      RECT  32.17 58.86 32.69 59.38 ;
      RECT  32.17 28.08 32.69 28.6 ;
      RECT  32.17 48.6 32.69 49.12 ;
      RECT  32.69 30.055 33.21 30.575 ;
      RECT  39.04 58.86 39.56 59.38 ;
      RECT  39.04 48.6 39.56 49.12 ;
      RECT  5.18 38.34 5.7 38.86 ;
      RECT  32.17 110.16 32.69 110.68 ;
      RECT  5.18 69.12 5.7 69.64 ;
      RECT  39.04 110.16 39.56 110.68 ;
      RECT  39.04 38.34 39.56 38.86 ;
      RECT  32.17 69.12 32.69 69.64 ;
      RECT  32.17 79.38 32.69 79.9 ;
      RECT  32.17 89.64 32.69 90.16 ;
      RECT  39.04 89.64 39.56 90.16 ;
      RECT  5.18 48.6 5.7 49.12 ;
      RECT  39.04 79.38 39.56 79.9 ;
      RECT  39.04 105.03 39.56 105.55 ;
      RECT  39.04 74.25 39.56 74.77 ;
      RECT  39.04 33.21 39.56 33.73 ;
      RECT  32.17 43.47 32.69 43.99 ;
      RECT  12.28 33.21 12.8 33.73 ;
      RECT  12.28 53.73 12.8 54.25 ;
      RECT  12.28 74.25 12.8 74.77 ;
      RECT  32.17 33.21 32.69 33.73 ;
      RECT  32.17 74.25 32.69 74.77 ;
      RECT  5.18 33.21 5.7 33.73 ;
      RECT  39.04 84.51 39.56 85.03 ;
      RECT  32.17 63.99 32.69 64.51 ;
      RECT  5.18 63.99 5.7 64.51 ;
      RECT  39.04 63.99 39.56 64.51 ;
      RECT  12.28 43.47 12.8 43.99 ;
      RECT  32.17 53.73 32.69 54.25 ;
      RECT  39.04 115.29 39.56 115.81 ;
      RECT  32.17 94.77 32.69 95.29 ;
      RECT  39.04 94.77 39.56 95.29 ;
      RECT  39.04 43.47 39.56 43.99 ;
      RECT  12.28 63.99 12.8 64.51 ;
      RECT  12.28 84.51 12.8 85.03 ;
      RECT  32.17 115.29 32.69 115.81 ;
      RECT  32.17 84.51 32.69 85.03 ;
      RECT  5.18 53.73 5.7 54.25 ;
      RECT  5.18 84.51 5.7 85.03 ;
      RECT  5.18 43.47 5.7 43.99 ;
      RECT  39.04 53.73 39.56 54.25 ;
      RECT  5.18 74.25 5.7 74.77 ;
      RECT  32.17 105.03 32.69 105.55 ;
      RECT  0.0 13.26 46.71 13.56 ;
      RECT  12.28 79.38 12.8 79.9 ;
      RECT  44.49 58.855 45.01 59.375 ;
      RECT  39.04 48.6 39.56 49.12 ;
      RECT  54.89 38.345 55.41 38.865 ;
      RECT  54.89 99.895 55.41 100.415 ;
      RECT  54.89 110.155 55.41 110.675 ;
      RECT  39.04 110.16 39.56 110.68 ;
      RECT  32.17 110.16 32.69 110.68 ;
      RECT  44.49 58.865 45.01 59.385 ;
      RECT  32.17 69.12 32.69 69.64 ;
      RECT  54.89 110.165 55.41 110.685 ;
      RECT  52.29 120.415 52.81 120.935 ;
      RECT  44.49 99.905 45.01 100.425 ;
      RECT  44.49 89.645 45.01 90.165 ;
      RECT  44.49 79.375 45.01 79.895 ;
      RECT  44.49 110.165 45.01 110.685 ;
      RECT  32.17 48.6 32.69 49.12 ;
      RECT  54.89 89.645 55.41 90.165 ;
      RECT  54.89 69.115 55.41 69.635 ;
      RECT  12.28 38.34 12.8 38.86 ;
      RECT  54.89 58.865 55.41 59.385 ;
      RECT  39.04 99.9 39.56 100.42 ;
      RECT  52.99 11.995 53.51 12.515 ;
      RECT  12.28 48.6 12.8 49.12 ;
      RECT  54.89 48.595 55.41 49.115 ;
      RECT  49.69 120.415 50.21 120.935 ;
      RECT  5.18 69.12 5.7 69.64 ;
      RECT  44.49 38.345 45.01 38.865 ;
      RECT  39.04 79.38 39.56 79.9 ;
      RECT  39.04 58.86 39.56 59.38 ;
      RECT  39.04 69.12 39.56 69.64 ;
      RECT  54.89 79.375 55.41 79.895 ;
      RECT  54.89 58.855 55.41 59.375 ;
      RECT  32.17 89.64 32.69 90.16 ;
      RECT  44.49 79.385 45.01 79.905 ;
      RECT  50.485 20.5 51.005 21.02 ;
      RECT  54.89 79.385 55.41 79.905 ;
      RECT  47.09 28.075 47.61 28.595 ;
      RECT  5.18 79.38 5.7 79.9 ;
      RECT  44.49 89.635 45.01 90.155 ;
      RECT  55.21 5.545 55.73 6.065 ;
      RECT  44.49 38.335 45.01 38.855 ;
      RECT  44.49 69.125 45.01 69.645 ;
      RECT  54.89 89.635 55.41 90.155 ;
      RECT  32.69 30.055 33.21 30.575 ;
      RECT  44.49 48.595 45.01 49.115 ;
      RECT  44.49 28.075 45.01 28.595 ;
      RECT  50.39 11.995 50.91 12.515 ;
      RECT  52.29 28.075 52.81 28.595 ;
      RECT  44.49 110.155 45.01 110.675 ;
      RECT  12.28 69.12 12.8 69.64 ;
      RECT  54.89 69.125 55.41 69.645 ;
      RECT  54.89 120.415 55.41 120.935 ;
      RECT  54.89 28.085 55.41 28.605 ;
      RECT  49.69 28.075 50.21 28.595 ;
      RECT  32.17 58.86 32.69 59.38 ;
      RECT  32.17 99.9 32.69 100.42 ;
      RECT  39.04 38.34 39.56 38.86 ;
      RECT  5.18 48.6 5.7 49.12 ;
      RECT  54.89 28.075 55.41 28.595 ;
      RECT  44.49 48.605 45.01 49.125 ;
      RECT  54.89 99.905 55.41 100.425 ;
      RECT  5.18 38.34 5.7 38.86 ;
      RECT  54.89 38.335 55.41 38.855 ;
      RECT  32.17 38.34 32.69 38.86 ;
      RECT  39.04 89.64 39.56 90.16 ;
      RECT  53.085 20.5 53.605 21.02 ;
      RECT  57.81 5.545 58.33 6.065 ;
      RECT  44.49 120.415 45.01 120.935 ;
      RECT  47.09 120.415 47.61 120.935 ;
      RECT  44.49 99.895 45.01 100.415 ;
      RECT  32.17 28.08 32.69 28.6 ;
      RECT  32.17 79.38 32.69 79.9 ;
      RECT  44.49 28.085 45.01 28.605 ;
      RECT  44.49 69.115 45.01 69.635 ;
      RECT  47.885 20.5 48.405 21.02 ;
      RECT  54.89 48.605 55.41 49.125 ;
      RECT  5.18 84.51 5.7 85.03 ;
      RECT  44.49 22.955 45.01 23.475 ;
      RECT  44.49 105.035 45.01 105.555 ;
      RECT  12.28 84.51 12.8 85.03 ;
      RECT  44.49 63.995 45.01 64.515 ;
      RECT  39.04 74.25 39.56 74.77 ;
      RECT  49.69 115.295 50.21 115.815 ;
      RECT  47.09 22.955 47.61 23.475 ;
      RECT  54.89 43.475 55.41 43.995 ;
      RECT  32.17 33.21 32.69 33.73 ;
      RECT  44.49 53.735 45.01 54.255 ;
      RECT  52.29 115.295 52.81 115.815 ;
      RECT  54.89 94.775 55.41 95.295 ;
      RECT  54.89 53.725 55.41 54.245 ;
      RECT  54.89 74.255 55.41 74.775 ;
      RECT  54.89 22.955 55.41 23.475 ;
      RECT  50.39 7.535 50.91 8.055 ;
      RECT  32.17 115.29 32.69 115.81 ;
      RECT  44.49 63.985 45.01 64.505 ;
      RECT  54.89 94.765 55.41 95.285 ;
      RECT  44.49 105.025 45.01 105.545 ;
      RECT  44.49 74.245 45.01 74.765 ;
      RECT  39.04 105.03 39.56 105.55 ;
      RECT  5.18 74.25 5.7 74.77 ;
      RECT  55.21 -0.265 55.73 0.255 ;
      RECT  12.28 53.73 12.8 54.25 ;
      RECT  12.28 74.25 12.8 74.77 ;
      RECT  54.89 115.295 55.41 115.815 ;
      RECT  39.04 43.47 39.56 43.99 ;
      RECT  39.04 33.21 39.56 33.73 ;
      RECT  47.09 115.295 47.61 115.815 ;
      RECT  44.49 94.765 45.01 95.285 ;
      RECT  44.49 84.515 45.01 85.035 ;
      RECT  39.04 53.73 39.56 54.25 ;
      RECT  44.49 43.475 45.01 43.995 ;
      RECT  54.89 63.985 55.41 64.505 ;
      RECT  54.89 33.205 55.41 33.725 ;
      RECT  44.49 74.255 45.01 74.775 ;
      RECT  32.17 84.51 32.69 85.03 ;
      RECT  32.17 43.47 32.69 43.99 ;
      RECT  52.99 7.535 53.51 8.055 ;
      RECT  5.18 43.47 5.7 43.99 ;
      RECT  44.49 33.205 45.01 33.725 ;
      RECT  57.09 116.38 57.61 116.9 ;
      RECT  44.49 115.295 45.01 115.815 ;
      RECT  42.29 116.38 42.81 116.9 ;
      RECT  12.28 63.99 12.8 64.51 ;
      RECT  57.09 24.04 57.61 24.56 ;
      RECT  32.17 94.77 32.69 95.29 ;
      RECT  39.04 63.99 39.56 64.51 ;
      RECT  54.89 63.995 55.41 64.515 ;
      RECT  52.29 22.955 52.81 23.475 ;
      RECT  54.89 43.465 55.41 43.985 ;
      RECT  44.49 33.215 45.01 33.735 ;
      RECT  54.89 105.025 55.41 105.545 ;
      RECT  32.17 74.25 32.69 74.77 ;
      RECT  5.18 53.73 5.7 54.25 ;
      RECT  44.49 43.465 45.01 43.985 ;
      RECT  32.17 63.99 32.69 64.51 ;
      RECT  5.18 33.21 5.7 33.73 ;
      RECT  44.49 53.725 45.01 54.245 ;
      RECT  39.04 115.29 39.56 115.81 ;
      RECT  54.89 53.735 55.41 54.255 ;
      RECT  39.04 84.51 39.56 85.03 ;
      RECT  42.29 24.04 42.81 24.56 ;
      RECT  44.49 94.775 45.01 95.295 ;
      RECT  54.89 84.505 55.41 85.025 ;
      RECT  44.49 84.505 45.01 85.025 ;
      RECT  57.81 -0.265 58.33 0.255 ;
      RECT  12.28 33.21 12.8 33.73 ;
      RECT  54.89 115.285 55.41 115.805 ;
      RECT  54.89 84.515 55.41 85.035 ;
      RECT  54.89 105.035 55.41 105.555 ;
      RECT  54.89 74.245 55.41 74.765 ;
      RECT  32.17 105.03 32.69 105.55 ;
      RECT  12.28 43.47 12.8 43.99 ;
      RECT  32.17 53.73 32.69 54.25 ;
      RECT  39.04 94.77 39.56 95.29 ;
      RECT  54.89 33.215 55.41 33.735 ;
      RECT  49.69 22.955 50.21 23.475 ;
      RECT  44.49 115.285 45.01 115.805 ;
      RECT  5.18 63.99 5.7 64.51 ;
      RECT  -55.65 -6.885 -55.13 -6.365 ;
      RECT  -55.65 -6.875 -55.13 -6.355 ;
      RECT  -55.71 -2.785 -55.19 -2.265 ;
      RECT  -55.71 -10.975 -55.19 -10.455 ;
      RECT  -45.17 31.35 -45.69 31.87 ;
      RECT  -45.17 81.75 -45.69 82.27 ;
      RECT  -45.17 81.75 -45.69 82.27 ;
      RECT  -51.45 98.55 -51.97 99.07 ;
      RECT  -45.17 64.95 -45.69 65.47 ;
      RECT  -45.17 48.15 -45.69 48.67 ;
      RECT  -51.45 48.15 -51.97 48.67 ;
      RECT  -45.17 98.55 -45.69 99.07 ;
      RECT  -51.45 31.35 -51.97 31.87 ;
      RECT  -45.17 31.35 -45.69 31.87 ;
      RECT  -51.45 81.75 -51.97 82.27 ;
      RECT  -51.45 81.75 -51.97 82.27 ;
      RECT  -51.45 64.95 -51.97 65.47 ;
      RECT  -51.45 31.35 -51.97 31.87 ;
      RECT  -45.17 73.35 -45.69 73.87 ;
      RECT  -51.45 73.35 -51.97 73.87 ;
      RECT  -45.17 39.75 -45.69 40.27 ;
      RECT  -51.45 56.55 -51.97 57.07 ;
      RECT  -51.45 39.75 -51.97 40.27 ;
      RECT  -51.45 90.15 -51.97 90.67 ;
      RECT  -45.17 22.95 -45.69 23.47 ;
      RECT  -45.17 56.55 -45.69 57.07 ;
      RECT  -51.45 22.95 -51.97 23.47 ;
      RECT  -45.17 90.15 -45.69 90.67 ;
      RECT  -51.97 31.35 -51.45 31.87 ;
      RECT  -51.97 98.55 -51.45 99.07 ;
      RECT  -55.65 -6.875 -55.13 -6.355 ;
      RECT  -51.97 64.95 -51.45 65.47 ;
      RECT  -45.69 31.35 -45.17 31.87 ;
      RECT  -45.69 98.55 -45.17 99.07 ;
      RECT  -45.69 64.95 -45.17 65.47 ;
      RECT  -45.69 81.75 -45.17 82.27 ;
      RECT  -55.65 -6.885 -55.13 -6.365 ;
      RECT  -51.97 48.15 -51.45 48.67 ;
      RECT  -45.69 48.15 -45.17 48.67 ;
      RECT  -51.97 81.75 -51.45 82.27 ;
      RECT  -51.97 73.35 -51.45 73.87 ;
      RECT  -45.69 73.35 -45.17 73.87 ;
      RECT  -51.97 90.15 -51.45 90.67 ;
      RECT  -51.97 22.95 -51.45 23.47 ;
      RECT  -51.97 39.75 -51.45 40.27 ;
      RECT  -45.69 90.15 -45.17 90.67 ;
      RECT  -55.71 -10.975 -55.19 -10.455 ;
      RECT  -45.69 22.95 -45.17 23.47 ;
      RECT  -45.69 39.75 -45.17 40.27 ;
      RECT  -55.71 -2.785 -55.19 -2.265 ;
      RECT  -51.97 56.55 -51.45 57.07 ;
      RECT  -45.69 56.55 -45.17 57.07 ;
      RECT  -14.03 101.8 -1.32 102.1 ;
      RECT  -7.905 112.025 -7.385 112.545 ;
      RECT  -7.905 112.015 -7.385 112.535 ;
      RECT  -7.905 103.845 -7.385 104.365 ;
      RECT  -7.905 103.835 -7.385 104.355 ;
      RECT  -8.025 107.935 -7.505 108.455 ;
      RECT  -8.025 107.925 -7.505 108.445 ;
      RECT  -8.025 99.745 -7.505 100.265 ;
      RECT  -8.025 116.115 -7.505 116.635 ;
      RECT  11.39 -8.92 36.81 -8.62 ;
      RECT  17.515 -6.885 18.035 -6.365 ;
      RECT  30.225 -6.885 30.745 -6.365 ;
      RECT  30.105 -10.975 30.625 -10.455 ;
      RECT  17.395 -10.975 17.915 -10.455 ;
   LAYER  m4 ;
   END
   END    sram_2_16_sky130A
END    LIBRARY
