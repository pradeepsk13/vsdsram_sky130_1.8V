magic
tech sky130A
timestamp 1606127284
<< nwell >>
rect 117 564 564 771
rect 748 564 1341 771
<< nmos >>
rect 185 217 200 259
rect 335 217 350 259
rect 481 217 496 259
rect 645 200 660 284
rect 816 217 831 259
rect 966 217 981 259
rect 1112 217 1127 259
rect 1276 185 1291 269
<< pmos >>
rect 185 584 200 639
rect 335 584 350 639
rect 481 584 496 639
rect 816 584 831 639
rect 966 584 981 639
rect 1112 584 1127 639
<< ndiff >>
rect 135 247 185 259
rect 135 230 150 247
rect 167 230 185 247
rect 135 217 185 230
rect 200 247 250 259
rect 200 230 218 247
rect 235 230 250 247
rect 200 217 250 230
rect 285 247 335 259
rect 285 230 300 247
rect 317 230 335 247
rect 285 217 335 230
rect 350 247 400 259
rect 350 230 368 247
rect 385 230 400 247
rect 350 217 400 230
rect 431 247 481 259
rect 431 230 446 247
rect 463 230 481 247
rect 431 217 481 230
rect 496 247 546 259
rect 496 230 514 247
rect 531 230 546 247
rect 496 217 546 230
rect 595 247 645 284
rect 595 230 610 247
rect 627 230 645 247
rect 595 200 645 230
rect 660 247 710 284
rect 660 230 678 247
rect 695 230 710 247
rect 660 200 710 230
rect 766 247 816 259
rect 766 230 781 247
rect 798 230 816 247
rect 766 217 816 230
rect 831 247 881 259
rect 831 230 849 247
rect 866 230 881 247
rect 831 217 881 230
rect 916 247 966 259
rect 916 230 931 247
rect 948 230 966 247
rect 916 217 966 230
rect 981 247 1020 259
rect 981 230 999 247
rect 1016 230 1020 247
rect 981 217 1020 230
rect 1065 247 1112 259
rect 1065 230 1077 247
rect 1094 230 1112 247
rect 1065 217 1112 230
rect 1127 247 1177 259
rect 1127 230 1145 247
rect 1162 230 1177 247
rect 1127 217 1177 230
rect 1226 247 1276 269
rect 1226 230 1241 247
rect 1258 230 1276 247
rect 1226 185 1276 230
rect 1291 247 1341 269
rect 1291 230 1309 247
rect 1326 230 1341 247
rect 1291 185 1341 230
<< pdiff >>
rect 135 620 185 639
rect 135 603 150 620
rect 167 603 185 620
rect 135 584 185 603
rect 200 620 250 639
rect 200 603 218 620
rect 235 603 250 620
rect 200 584 250 603
rect 285 620 335 639
rect 285 603 300 620
rect 317 603 335 620
rect 285 584 335 603
rect 350 620 400 639
rect 350 603 368 620
rect 385 603 400 620
rect 350 584 400 603
rect 431 620 481 639
rect 431 603 446 620
rect 463 603 481 620
rect 431 584 481 603
rect 496 620 546 639
rect 496 603 514 620
rect 531 603 546 620
rect 496 584 546 603
rect 766 620 816 639
rect 766 603 781 620
rect 798 603 816 620
rect 766 584 816 603
rect 831 620 881 639
rect 831 603 849 620
rect 866 603 881 620
rect 831 584 881 603
rect 916 620 966 639
rect 916 603 931 620
rect 948 603 966 620
rect 916 584 966 603
rect 981 620 1031 639
rect 981 603 999 620
rect 1016 603 1031 620
rect 981 584 1031 603
rect 1062 620 1112 639
rect 1062 603 1077 620
rect 1094 603 1112 620
rect 1062 584 1112 603
rect 1127 620 1177 639
rect 1127 603 1145 620
rect 1162 603 1177 620
rect 1127 584 1177 603
<< ndiffc >>
rect 150 230 167 247
rect 218 230 235 247
rect 300 230 317 247
rect 368 230 385 247
rect 446 230 463 247
rect 514 230 531 247
rect 610 230 627 247
rect 678 230 695 247
rect 781 230 798 247
rect 849 230 866 247
rect 931 230 948 247
rect 999 230 1016 247
rect 1077 230 1094 247
rect 1145 230 1162 247
rect 1241 230 1258 247
rect 1309 230 1326 247
<< pdiffc >>
rect 150 603 167 620
rect 218 603 235 620
rect 300 603 317 620
rect 368 603 385 620
rect 446 603 463 620
rect 514 603 531 620
rect 781 603 798 620
rect 849 603 866 620
rect 931 603 948 620
rect 999 603 1016 620
rect 1077 603 1094 620
rect 1145 603 1162 620
<< psubdiff >>
rect 173 144 214 156
rect 173 127 185 144
rect 202 127 214 144
rect 173 115 214 127
rect 323 144 364 156
rect 323 127 335 144
rect 352 127 364 144
rect 323 115 364 127
rect 469 144 510 156
rect 469 127 481 144
rect 498 127 510 144
rect 469 115 510 127
rect 633 144 674 156
rect 633 127 645 144
rect 662 127 674 144
rect 633 115 674 127
rect 804 144 845 156
rect 804 127 816 144
rect 833 127 845 144
rect 804 115 845 127
rect 954 144 995 156
rect 954 127 966 144
rect 983 127 995 144
rect 954 115 995 127
rect 1100 144 1141 156
rect 1100 127 1112 144
rect 1129 127 1141 144
rect 1100 115 1141 127
rect 1264 144 1305 156
rect 1264 127 1276 144
rect 1293 127 1305 144
rect 1264 115 1305 127
<< nsubdiff >>
rect 160 726 213 744
rect 160 709 178 726
rect 195 709 213 726
rect 160 691 213 709
rect 310 726 363 744
rect 310 709 328 726
rect 345 709 363 726
rect 310 691 363 709
rect 456 726 509 744
rect 456 709 474 726
rect 491 709 509 726
rect 456 691 509 709
rect 791 726 844 744
rect 791 709 809 726
rect 826 709 844 726
rect 791 691 844 709
rect 941 726 994 744
rect 941 709 959 726
rect 976 709 994 726
rect 941 691 994 709
rect 1087 726 1140 744
rect 1087 709 1105 726
rect 1122 709 1140 726
rect 1087 691 1140 709
rect 1225 726 1278 744
rect 1225 709 1243 726
rect 1260 709 1278 726
rect 1225 691 1278 709
<< psubdiffcont >>
rect 185 127 202 144
rect 335 127 352 144
rect 481 127 498 144
rect 645 127 662 144
rect 816 127 833 144
rect 966 127 983 144
rect 1112 127 1129 144
rect 1276 127 1293 144
<< nsubdiffcont >>
rect 178 709 195 726
rect 328 709 345 726
rect 474 709 491 726
rect 809 709 826 726
rect 959 709 976 726
rect 1105 709 1122 726
rect 1243 709 1260 726
<< poly >>
rect 185 639 200 654
rect 335 639 350 654
rect 481 639 496 654
rect 816 639 831 654
rect 966 639 981 654
rect 1112 639 1127 654
rect 127 327 160 335
rect 127 310 135 327
rect 152 325 160 327
rect 185 325 200 584
rect 335 520 350 584
rect 326 512 359 520
rect 326 495 334 512
rect 351 495 359 512
rect 326 487 359 495
rect 152 310 200 325
rect 127 302 160 310
rect 185 259 200 310
rect 335 259 350 487
rect 481 388 496 584
rect 758 511 791 519
rect 758 494 766 511
rect 783 509 791 511
rect 816 509 831 584
rect 966 520 981 584
rect 783 494 831 509
rect 758 486 791 494
rect 471 380 504 388
rect 471 363 479 380
rect 496 363 504 380
rect 471 355 504 363
rect 481 259 496 355
rect 577 327 610 335
rect 577 310 585 327
rect 602 325 610 327
rect 602 310 660 325
rect 577 302 610 310
rect 645 284 660 310
rect 185 202 200 217
rect 335 202 350 217
rect 481 202 496 217
rect 816 259 831 494
rect 957 512 990 520
rect 957 495 965 512
rect 982 495 990 512
rect 957 487 990 495
rect 966 259 981 487
rect 1112 401 1127 584
rect 1094 393 1127 401
rect 1094 376 1102 393
rect 1119 376 1127 393
rect 1094 368 1127 376
rect 1112 259 1127 368
rect 1208 327 1241 335
rect 1208 310 1216 327
rect 1233 325 1241 327
rect 1233 310 1291 325
rect 1208 302 1241 310
rect 1276 269 1291 310
rect 816 202 831 217
rect 966 202 981 217
rect 1112 202 1127 217
rect 645 185 660 200
rect 1276 170 1291 185
<< polycont >>
rect 135 310 152 327
rect 334 495 351 512
rect 766 494 783 511
rect 479 363 496 380
rect 585 310 602 327
rect 965 495 982 512
rect 1102 376 1119 393
rect 1216 310 1233 327
<< locali >>
rect 117 727 1341 739
rect 117 726 610 727
rect 117 709 178 726
rect 195 709 235 726
rect 252 709 328 726
rect 345 709 385 726
rect 402 709 474 726
rect 491 709 531 726
rect 548 710 610 726
rect 627 710 669 727
rect 686 710 717 727
rect 734 726 1341 727
rect 734 710 809 726
rect 548 709 809 710
rect 826 709 866 726
rect 883 709 959 726
rect 976 709 1016 726
rect 1033 709 1105 726
rect 1122 709 1162 726
rect 1179 709 1243 726
rect 1260 709 1300 726
rect 1317 709 1341 726
rect 117 694 1341 709
rect 150 639 170 694
rect 300 639 320 694
rect 781 639 801 694
rect 931 639 951 694
rect 142 620 175 639
rect 142 603 150 620
rect 167 603 175 620
rect 142 595 175 603
rect 210 620 243 639
rect 210 603 218 620
rect 235 603 243 620
rect 210 595 243 603
rect 292 620 325 639
rect 292 603 300 620
rect 317 603 325 620
rect 292 595 325 603
rect 360 620 471 639
rect 360 603 368 620
rect 385 603 446 620
rect 463 603 471 620
rect 360 595 471 603
rect 506 620 539 639
rect 506 603 514 620
rect 531 603 539 620
rect 506 595 539 603
rect 773 620 806 639
rect 773 603 781 620
rect 798 603 806 620
rect 773 595 806 603
rect 841 620 874 639
rect 841 603 849 620
rect 866 603 874 620
rect 841 595 874 603
rect 923 620 956 639
rect 923 603 931 620
rect 948 603 956 620
rect 923 595 956 603
rect 991 620 1102 639
rect 991 603 999 620
rect 1016 603 1077 620
rect 1094 603 1102 620
rect 991 595 1102 603
rect 1137 620 1170 639
rect 1137 603 1145 620
rect 1162 603 1170 620
rect 1137 595 1170 603
rect 215 513 235 595
rect 515 570 535 595
rect 508 564 538 570
rect 508 547 515 564
rect 532 547 538 564
rect 508 541 538 547
rect 326 513 359 520
rect 758 513 791 519
rect 215 512 791 513
rect 215 495 334 512
rect 351 511 791 512
rect 351 495 766 511
rect 215 494 766 495
rect 783 494 791 511
rect 215 493 791 494
rect 47 327 77 332
rect 127 327 160 335
rect 47 325 135 327
rect 47 308 54 325
rect 71 310 135 325
rect 152 310 160 327
rect 71 308 160 310
rect 47 307 160 308
rect 47 302 77 307
rect 127 302 160 307
rect 215 255 235 493
rect 326 487 359 493
rect 758 486 791 493
rect 846 513 866 595
rect 1146 570 1166 595
rect 1139 564 1169 570
rect 1139 547 1146 564
rect 1163 547 1169 564
rect 1139 541 1169 547
rect 957 513 990 520
rect 846 512 990 513
rect 846 495 965 512
rect 982 495 990 512
rect 846 493 990 495
rect 678 464 708 470
rect 678 447 685 464
rect 702 447 708 464
rect 678 441 708 447
rect 633 391 663 397
rect 471 385 504 388
rect 633 385 640 391
rect 277 380 307 385
rect 471 380 640 385
rect 277 378 479 380
rect 277 361 284 378
rect 301 363 479 378
rect 496 374 640 380
rect 657 374 663 391
rect 496 368 663 374
rect 496 363 504 368
rect 301 361 504 363
rect 277 360 504 361
rect 277 355 307 360
rect 471 355 504 360
rect 508 331 538 337
rect 508 330 515 331
rect 375 314 515 330
rect 532 330 538 331
rect 577 330 610 335
rect 532 327 610 330
rect 532 314 585 327
rect 375 310 585 314
rect 602 310 610 327
rect 375 255 395 310
rect 508 308 538 310
rect 515 255 535 308
rect 577 302 610 310
rect 680 255 700 441
rect 846 255 866 493
rect 957 487 990 493
rect 1031 465 1061 470
rect 1294 465 1324 470
rect 1031 464 1324 465
rect 1031 447 1038 464
rect 1055 447 1301 464
rect 1318 447 1324 464
rect 1031 445 1324 447
rect 1031 441 1061 445
rect 1294 441 1324 445
rect 1094 393 1127 401
rect 1094 376 1102 393
rect 1119 376 1127 393
rect 1094 368 1127 376
rect 1139 331 1169 337
rect 1139 330 1146 331
rect 995 314 1146 330
rect 1163 330 1169 331
rect 1208 330 1241 335
rect 1163 327 1241 330
rect 1163 314 1216 327
rect 995 310 1216 314
rect 1233 310 1241 327
rect 995 255 1015 310
rect 1139 308 1169 310
rect 1145 255 1165 308
rect 1208 302 1241 310
rect 1310 327 1340 333
rect 1310 310 1317 327
rect 1334 310 1340 327
rect 1310 304 1340 310
rect 1310 255 1330 304
rect 142 247 175 255
rect 142 230 150 247
rect 167 230 175 247
rect 142 217 175 230
rect 210 247 243 255
rect 210 230 218 247
rect 235 230 243 247
rect 210 217 243 230
rect 292 247 325 255
rect 292 230 300 247
rect 317 230 325 247
rect 292 217 325 230
rect 360 247 400 255
rect 360 230 368 247
rect 385 230 400 247
rect 360 217 400 230
rect 431 247 471 255
rect 431 230 446 247
rect 463 230 471 247
rect 431 217 471 230
rect 506 247 539 255
rect 506 230 514 247
rect 531 230 539 247
rect 506 217 539 230
rect 602 247 635 255
rect 602 230 610 247
rect 627 230 635 247
rect 602 217 635 230
rect 670 247 703 255
rect 670 230 678 247
rect 695 230 703 247
rect 670 217 703 230
rect 773 247 806 255
rect 773 230 781 247
rect 798 230 806 247
rect 773 217 806 230
rect 841 247 874 255
rect 841 230 849 247
rect 866 230 874 247
rect 841 217 874 230
rect 923 247 956 255
rect 923 230 931 247
rect 948 230 956 247
rect 923 217 956 230
rect 991 247 1020 255
rect 991 230 999 247
rect 1016 230 1020 247
rect 991 217 1020 230
rect 1065 247 1102 255
rect 1065 230 1077 247
rect 1094 230 1102 247
rect 1065 217 1102 230
rect 1137 247 1170 255
rect 1137 230 1145 247
rect 1162 230 1170 247
rect 1137 217 1170 230
rect 1233 247 1266 255
rect 1233 230 1241 247
rect 1258 230 1266 247
rect 1233 217 1266 230
rect 1301 247 1334 255
rect 1301 230 1309 247
rect 1326 230 1334 247
rect 1301 217 1334 230
rect 145 152 165 217
rect 300 152 320 217
rect 440 152 460 217
rect 610 152 630 217
rect 776 152 796 217
rect 931 152 951 217
rect 1070 152 1090 217
rect 1241 152 1261 217
rect 117 144 1341 152
rect 117 127 150 144
rect 167 127 185 144
rect 202 127 228 144
rect 245 127 300 144
rect 317 127 335 144
rect 352 127 378 144
rect 395 127 446 144
rect 463 127 481 144
rect 498 127 524 144
rect 541 127 610 144
rect 627 127 645 144
rect 662 127 688 144
rect 705 127 781 144
rect 798 127 816 144
rect 833 127 859 144
rect 876 127 931 144
rect 948 127 966 144
rect 983 127 1009 144
rect 1026 127 1077 144
rect 1094 127 1112 144
rect 1129 127 1155 144
rect 1172 127 1241 144
rect 1258 127 1276 144
rect 1293 127 1319 144
rect 1336 127 1341 144
rect 117 119 1341 127
<< viali >>
rect 235 709 252 726
rect 385 709 402 726
rect 531 709 548 726
rect 610 710 627 727
rect 669 710 686 727
rect 717 710 734 727
rect 866 709 883 726
rect 1016 709 1033 726
rect 1162 709 1179 726
rect 1300 709 1317 726
rect 515 547 532 564
rect 54 308 71 325
rect 1146 547 1163 564
rect 685 447 702 464
rect 284 361 301 378
rect 640 374 657 391
rect 515 314 532 331
rect 1038 447 1055 464
rect 1301 447 1318 464
rect 1102 376 1119 393
rect 1146 314 1163 331
rect 1317 310 1334 327
rect 150 127 167 144
rect 228 127 245 144
rect 300 127 317 144
rect 378 127 395 144
rect 446 127 463 144
rect 524 127 541 144
rect 610 127 627 144
rect 688 127 705 144
rect 781 127 798 144
rect 859 127 876 144
rect 931 127 948 144
rect 1009 127 1026 144
rect 1077 127 1094 144
rect 1155 127 1172 144
rect 1241 127 1258 144
rect 1319 127 1336 144
<< metal1 >>
rect 117 727 1341 739
rect 117 726 610 727
rect 117 709 235 726
rect 252 709 385 726
rect 402 709 531 726
rect 548 710 610 726
rect 627 710 669 727
rect 686 710 717 727
rect 734 726 1341 727
rect 734 710 866 726
rect 548 709 866 710
rect 883 709 1016 726
rect 1033 709 1162 726
rect 1179 709 1300 726
rect 1317 709 1341 726
rect 117 694 1341 709
rect 508 564 538 570
rect 508 547 515 564
rect 532 547 538 564
rect 277 380 307 385
rect 104 378 307 380
rect 104 361 284 378
rect 301 361 307 378
rect 104 360 307 361
rect 277 355 307 360
rect 47 325 77 332
rect 47 308 54 325
rect 71 308 77 325
rect 508 331 538 547
rect 1139 564 1169 570
rect 1139 547 1146 564
rect 1163 547 1169 564
rect 1139 541 1169 547
rect 678 464 1061 470
rect 678 447 685 464
rect 702 447 1038 464
rect 1055 447 1061 464
rect 678 441 1061 447
rect 1094 397 1127 401
rect 633 393 1127 397
rect 633 391 1102 393
rect 633 374 640 391
rect 657 376 1102 391
rect 1119 376 1127 393
rect 657 374 1127 376
rect 633 368 1127 374
rect 1143 337 1169 541
rect 1294 464 1324 470
rect 1294 447 1301 464
rect 1318 447 1324 464
rect 1294 441 1324 447
rect 508 314 515 331
rect 532 314 538 331
rect 508 308 538 314
rect 1139 331 1169 337
rect 1139 314 1146 331
rect 1163 314 1169 331
rect 1139 308 1169 314
rect 1310 327 1340 333
rect 1310 310 1317 327
rect 1334 310 1340 327
rect 47 302 77 308
rect 1310 304 1340 310
rect 117 144 1341 152
rect 117 127 150 144
rect 167 127 228 144
rect 245 127 300 144
rect 317 127 378 144
rect 395 127 446 144
rect 463 127 524 144
rect 541 127 610 144
rect 627 127 688 144
rect 705 127 781 144
rect 798 127 859 144
rect 876 127 931 144
rect 948 127 1009 144
rect 1026 127 1077 144
rect 1094 127 1155 144
rect 1172 127 1241 144
rect 1258 127 1319 144
rect 1336 127 1341 144
rect 117 119 1341 127
<< labels >>
flabel locali s 1304 451 1314 460 0 FreeSans 600 0 0 0 blb
port 0 nsew
flabel locali s 1321 315 1331 324 0 FreeSans 600 0 0 0 bl
port 1 nsew
flabel metal1 s 552 124 591 143 0 FreeSans 400 0 0 0 gnd
port 2 nsew
flabel metal1 s 569 714 608 733 0 FreeSans 400 0 0 0 vdd
port 3 nsew
flabel locali s 136 311 146 322 0 FreeSans 400 0 0 0 din
port 4 nsew
flabel locali s 482 368 492 379 0 FreeSans 400 0 0 0 wb
port 5 nsew
flabel locali s 223 440 233 451 0 FreeSans 200 0 0 0 net1
flabel locali s 871 499 881 510 0 FreeSans 200 0 0 0 net3
flabel locali s 1149 318 1159 329 0 FreeSans 200 0 0 0 net4
flabel locali s 517 316 527 327 0 FreeSans 200 0 0 0 net2
flabel locali s 406 606 416 617 0 FreeSans 200 0 0 0 net5
flabel locali s 1038 606 1048 617 0 FreeSans 200 0 0 0 net6
<< end >>
