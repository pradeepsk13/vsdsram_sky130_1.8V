magic
tech sky130A
timestamp 1606126701
<< nwell >>
rect -10 285 78 292
rect 1126 289 1309 291
rect 877 288 1309 289
rect 566 287 1309 288
rect 441 286 1309 287
rect 345 285 1309 286
rect -10 217 1309 285
rect -10 185 1310 217
rect -8 113 1310 185
rect 440 112 1310 113
rect 566 110 1309 112
rect -8 -247 346 -76
<< nmos >>
rect 45 20 60 62
rect 160 20 175 62
rect 275 20 290 62
rect 390 -22 405 62
rect 687 -85 702 41
rect 800 -84 815 42
rect 1230 19 1245 61
rect 1040 -86 1055 14
rect 800 -210 815 -168
rect 952 -186 967 -144
rect 1092 -185 1107 -143
rect 686 -263 701 -221
rect 45 -381 60 -339
rect 160 -381 175 -339
rect 275 -381 290 -339
rect 390 -423 405 -339
<< pmos >>
rect 45 131 60 186
rect 160 131 175 186
rect 275 131 290 186
rect 390 148 405 203
rect 505 148 520 203
rect 687 131 702 186
rect 800 131 815 186
rect 958 131 973 186
rect 1071 131 1086 231
rect 1230 130 1245 185
rect 45 -229 60 -174
rect 160 -229 175 -174
rect 275 -229 290 -174
<< ndiff >>
rect 10 47 45 62
rect 10 30 18 47
rect 35 30 45 47
rect 10 20 45 30
rect 60 47 95 62
rect 60 30 70 47
rect 87 30 95 47
rect 60 20 95 30
rect 125 47 160 62
rect 125 30 133 47
rect 150 30 160 47
rect 125 20 160 30
rect 175 47 210 62
rect 175 30 185 47
rect 202 30 210 47
rect 175 20 210 30
rect 240 47 275 62
rect 240 30 248 47
rect 265 30 275 47
rect 240 20 275 30
rect 290 47 325 62
rect 290 30 300 47
rect 317 30 325 47
rect 290 20 325 30
rect 355 47 390 62
rect 355 30 363 47
rect 380 30 390 47
rect 355 -22 390 30
rect 405 47 440 62
rect 405 30 415 47
rect 432 30 440 47
rect 405 -22 440 30
rect 652 26 687 41
rect 652 9 660 26
rect 677 9 687 26
rect 652 -85 687 9
rect 702 26 737 41
rect 702 9 712 26
rect 729 9 737 26
rect 702 -85 737 9
rect 765 27 800 42
rect 765 10 773 27
rect 790 10 800 27
rect 765 -84 800 10
rect 815 27 850 42
rect 1195 46 1230 61
rect 815 10 825 27
rect 842 10 850 27
rect 1195 29 1203 46
rect 1220 29 1230 46
rect 1195 19 1230 29
rect 1245 46 1280 61
rect 1245 29 1255 46
rect 1272 29 1280 46
rect 1245 19 1280 29
rect 815 -84 850 10
rect 1005 -59 1040 14
rect 1005 -76 1013 -59
rect 1030 -76 1040 -59
rect 1005 -86 1040 -76
rect 1055 -59 1090 14
rect 1055 -76 1065 -59
rect 1082 -76 1090 -59
rect 1055 -86 1090 -76
rect 917 -159 952 -144
rect 765 -183 800 -168
rect 765 -200 773 -183
rect 790 -200 800 -183
rect 765 -210 800 -200
rect 815 -183 850 -168
rect 815 -200 825 -183
rect 842 -200 850 -183
rect 917 -176 925 -159
rect 942 -176 952 -159
rect 917 -186 952 -176
rect 967 -159 1002 -144
rect 967 -176 977 -159
rect 994 -176 1002 -159
rect 967 -186 1002 -176
rect 1057 -158 1092 -143
rect 1057 -175 1065 -158
rect 1082 -175 1092 -158
rect 1057 -185 1092 -175
rect 1107 -158 1142 -143
rect 1107 -175 1117 -158
rect 1134 -175 1142 -158
rect 1107 -185 1142 -175
rect 815 -210 850 -200
rect 651 -236 686 -221
rect 651 -253 659 -236
rect 676 -253 686 -236
rect 651 -263 686 -253
rect 701 -236 736 -221
rect 701 -253 711 -236
rect 728 -253 736 -236
rect 701 -263 736 -253
rect 10 -354 45 -339
rect 10 -371 18 -354
rect 35 -371 45 -354
rect 10 -381 45 -371
rect 60 -354 95 -339
rect 60 -371 70 -354
rect 87 -371 95 -354
rect 60 -381 95 -371
rect 125 -354 160 -339
rect 125 -371 133 -354
rect 150 -371 160 -354
rect 125 -381 160 -371
rect 175 -354 210 -339
rect 175 -371 185 -354
rect 202 -371 210 -354
rect 175 -381 210 -371
rect 240 -354 275 -339
rect 240 -371 248 -354
rect 265 -371 275 -354
rect 240 -381 275 -371
rect 290 -354 325 -339
rect 290 -371 300 -354
rect 317 -371 325 -354
rect 290 -381 325 -371
rect 355 -354 390 -339
rect 355 -371 363 -354
rect 380 -371 390 -354
rect 355 -423 390 -371
rect 405 -354 440 -339
rect 405 -371 415 -354
rect 432 -371 440 -354
rect 405 -423 440 -371
<< pdiff >>
rect 10 164 45 186
rect 10 147 18 164
rect 35 147 45 164
rect 10 131 45 147
rect 60 164 95 186
rect 60 147 70 164
rect 87 147 95 164
rect 60 131 95 147
rect 125 164 160 186
rect 125 147 133 164
rect 150 147 160 164
rect 125 131 160 147
rect 175 164 210 186
rect 175 147 185 164
rect 202 147 210 164
rect 175 131 210 147
rect 240 164 275 186
rect 240 147 248 164
rect 265 147 275 164
rect 240 131 275 147
rect 290 164 325 186
rect 290 147 300 164
rect 317 147 325 164
rect 355 181 390 203
rect 355 164 363 181
rect 380 164 390 181
rect 355 148 390 164
rect 405 181 440 203
rect 405 164 415 181
rect 432 164 440 181
rect 405 148 440 164
rect 470 181 505 203
rect 470 164 478 181
rect 495 164 505 181
rect 470 148 505 164
rect 520 181 555 203
rect 1036 186 1071 231
rect 520 164 530 181
rect 547 164 555 181
rect 520 148 555 164
rect 652 164 687 186
rect 290 131 325 147
rect 652 147 660 164
rect 677 147 687 164
rect 652 131 687 147
rect 702 164 737 186
rect 702 147 712 164
rect 729 147 737 164
rect 702 131 737 147
rect 765 164 800 186
rect 765 147 773 164
rect 790 147 800 164
rect 765 131 800 147
rect 815 164 850 186
rect 815 147 825 164
rect 842 147 850 164
rect 815 131 850 147
rect 923 164 958 186
rect 923 147 931 164
rect 948 147 958 164
rect 923 131 958 147
rect 973 164 1071 186
rect 973 147 983 164
rect 1000 147 1044 164
rect 1061 147 1071 164
rect 973 131 1071 147
rect 1086 164 1121 231
rect 1086 147 1096 164
rect 1113 147 1121 164
rect 1086 131 1121 147
rect 1195 163 1230 185
rect 1195 146 1203 163
rect 1220 146 1230 163
rect 1195 130 1230 146
rect 1245 163 1280 185
rect 1245 146 1255 163
rect 1272 146 1280 163
rect 1245 130 1280 146
rect 10 -196 45 -174
rect 10 -213 18 -196
rect 35 -213 45 -196
rect 10 -229 45 -213
rect 60 -196 95 -174
rect 60 -213 70 -196
rect 87 -213 95 -196
rect 60 -229 95 -213
rect 125 -196 160 -174
rect 125 -213 133 -196
rect 150 -213 160 -196
rect 125 -229 160 -213
rect 175 -196 210 -174
rect 175 -213 185 -196
rect 202 -213 210 -196
rect 175 -229 210 -213
rect 240 -196 275 -174
rect 240 -213 248 -196
rect 265 -213 275 -196
rect 240 -229 275 -213
rect 290 -196 325 -174
rect 290 -213 300 -196
rect 317 -213 325 -196
rect 290 -229 325 -213
<< ndiffc >>
rect 18 30 35 47
rect 70 30 87 47
rect 133 30 150 47
rect 185 30 202 47
rect 248 30 265 47
rect 300 30 317 47
rect 363 30 380 47
rect 415 30 432 47
rect 660 9 677 26
rect 712 9 729 26
rect 773 10 790 27
rect 825 10 842 27
rect 1203 29 1220 46
rect 1255 29 1272 46
rect 1013 -76 1030 -59
rect 1065 -76 1082 -59
rect 773 -200 790 -183
rect 825 -200 842 -183
rect 925 -176 942 -159
rect 977 -176 994 -159
rect 1065 -175 1082 -158
rect 1117 -175 1134 -158
rect 659 -253 676 -236
rect 711 -253 728 -236
rect 18 -371 35 -354
rect 70 -371 87 -354
rect 133 -371 150 -354
rect 185 -371 202 -354
rect 248 -371 265 -354
rect 300 -371 317 -354
rect 363 -371 380 -354
rect 415 -371 432 -354
<< pdiffc >>
rect 18 147 35 164
rect 70 147 87 164
rect 133 147 150 164
rect 185 147 202 164
rect 248 147 265 164
rect 300 147 317 164
rect 363 164 380 181
rect 415 164 432 181
rect 478 164 495 181
rect 530 164 547 181
rect 660 147 677 164
rect 712 147 729 164
rect 773 147 790 164
rect 825 147 842 164
rect 931 147 948 164
rect 983 147 1000 164
rect 1044 147 1061 164
rect 1096 147 1113 164
rect 1203 146 1220 163
rect 1255 146 1272 163
rect 18 -213 35 -196
rect 70 -213 87 -196
rect 133 -213 150 -196
rect 185 -213 202 -196
rect 248 -213 265 -196
rect 300 -213 317 -196
<< psubdiff >>
rect 93 -25 134 -13
rect 93 -42 105 -25
rect 122 -42 134 -25
rect 93 -54 134 -42
rect 210 -25 251 -13
rect 210 -42 222 -25
rect 239 -42 251 -25
rect 210 -54 251 -42
rect 486 -25 527 -13
rect 486 -42 498 -25
rect 515 -42 527 -25
rect 486 -54 527 -42
rect 1271 -23 1312 -11
rect 1271 -40 1283 -23
rect 1300 -40 1312 -23
rect 1271 -52 1312 -40
rect 90 -423 131 -411
rect 90 -440 102 -423
rect 119 -440 131 -423
rect 90 -452 131 -440
rect 245 -423 286 -411
rect 245 -440 257 -423
rect 274 -440 286 -423
rect 245 -452 286 -440
<< nsubdiff >>
rect 86 249 139 267
rect 86 232 104 249
rect 121 232 139 249
rect 86 215 139 232
rect 266 249 319 267
rect 266 232 284 249
rect 301 232 319 249
rect 266 215 319 232
rect 678 249 731 267
rect 678 232 696 249
rect 713 232 731 249
rect 678 215 731 232
rect 791 249 844 267
rect 791 232 809 249
rect 826 232 844 249
rect 791 215 844 232
rect 888 249 941 267
rect 888 232 906 249
rect 923 232 941 249
rect 888 215 941 232
rect 1174 249 1227 267
rect 1174 232 1192 249
rect 1209 232 1227 249
rect 1174 215 1227 232
rect 87 -112 140 -94
rect 87 -129 105 -112
rect 122 -129 140 -112
rect 87 -146 140 -129
rect 200 -112 253 -94
rect 200 -129 218 -112
rect 235 -129 253 -112
rect 200 -146 253 -129
<< psubdiffcont >>
rect 105 -42 122 -25
rect 222 -42 239 -25
rect 498 -42 515 -25
rect 1283 -40 1300 -23
rect 102 -440 119 -423
rect 257 -440 274 -423
<< nsubdiffcont >>
rect 104 232 121 249
rect 284 232 301 249
rect 696 232 713 249
rect 809 232 826 249
rect 906 232 923 249
rect 1192 232 1209 249
rect 105 -129 122 -112
rect 218 -129 235 -112
<< poly >>
rect 390 215 520 230
rect 958 250 1086 265
rect 390 203 405 215
rect 505 203 520 215
rect 45 186 60 200
rect 160 186 175 200
rect 275 186 290 200
rect 687 186 702 200
rect 800 186 815 200
rect 958 186 973 250
rect 1071 231 1086 250
rect -111 100 -78 108
rect -111 83 -103 100
rect -86 95 -78 100
rect 45 95 60 131
rect -86 83 60 95
rect -111 80 60 83
rect -111 75 -78 80
rect 45 62 60 80
rect 103 98 136 106
rect 103 81 111 98
rect 128 95 136 98
rect 160 95 175 131
rect 128 81 175 95
rect 103 80 175 81
rect 103 73 136 80
rect 160 62 175 80
rect 275 62 290 131
rect 390 129 405 148
rect 372 100 405 108
rect 505 107 520 148
rect 1230 185 1245 205
rect 372 83 380 100
rect 397 83 405 100
rect 372 75 405 83
rect 390 62 405 75
rect 496 99 529 107
rect 496 82 504 99
rect 521 82 529 99
rect 687 85 702 131
rect 800 115 815 131
rect 496 74 529 82
rect 654 77 702 85
rect 767 107 815 115
rect 767 90 775 107
rect 792 90 815 107
rect 767 82 815 90
rect 45 5 60 20
rect 160 -70 175 20
rect 45 -85 175 -70
rect 45 -174 60 -85
rect 160 -174 175 -160
rect 275 -174 290 20
rect 654 60 662 77
rect 679 60 702 77
rect 654 52 702 60
rect 687 41 702 52
rect 800 42 815 82
rect 958 105 973 131
rect 1071 106 1086 131
rect 958 97 991 105
rect 958 80 966 97
rect 983 80 991 97
rect 958 72 991 80
rect 1144 95 1177 103
rect 1144 78 1152 95
rect 1169 94 1177 95
rect 1230 94 1245 130
rect 1169 79 1245 94
rect 1169 78 1177 79
rect 1144 70 1177 78
rect 1032 56 1065 64
rect 1230 61 1245 79
rect 390 -40 405 -22
rect 1032 39 1040 56
rect 1057 39 1065 56
rect 1032 31 1065 39
rect 1040 14 1055 31
rect 687 -101 702 -85
rect 800 -101 815 -84
rect 1230 2 1245 19
rect 1040 -105 1055 -86
rect 952 -144 967 -128
rect 1092 -143 1107 -127
rect 800 -168 815 -152
rect 686 -221 701 -183
rect 45 -339 60 -229
rect 160 -266 175 -229
rect 275 -246 290 -229
rect 127 -274 175 -266
rect 127 -291 135 -274
rect 152 -291 175 -274
rect 257 -254 290 -246
rect 257 -271 265 -254
rect 282 -271 290 -254
rect 257 -279 290 -271
rect 127 -299 175 -291
rect 160 -339 175 -299
rect 275 -339 290 -279
rect 686 -280 701 -263
rect 800 -270 815 -210
rect 952 -213 967 -186
rect 1092 -204 1107 -185
rect 1083 -212 1116 -204
rect 943 -221 976 -213
rect 943 -238 951 -221
rect 968 -238 976 -221
rect 1083 -229 1091 -212
rect 1108 -229 1116 -212
rect 1083 -237 1116 -229
rect 943 -246 976 -238
rect 790 -278 823 -270
rect 790 -280 798 -278
rect 372 -299 405 -291
rect 686 -295 798 -280
rect 815 -295 823 -278
rect 372 -316 380 -299
rect 397 -316 405 -299
rect 790 -303 823 -295
rect 372 -324 405 -316
rect 390 -339 405 -324
rect 45 -396 60 -381
rect 160 -396 175 -381
rect 275 -396 290 -381
rect 390 -439 405 -423
<< polycont >>
rect -103 83 -86 100
rect 111 81 128 98
rect 380 83 397 100
rect 504 82 521 99
rect 775 90 792 107
rect 662 60 679 77
rect 966 80 983 97
rect 1152 78 1169 95
rect 1040 39 1057 56
rect 135 -291 152 -274
rect 265 -271 282 -254
rect 951 -238 968 -221
rect 1091 -229 1108 -212
rect 798 -295 815 -278
rect 380 -316 397 -299
<< locali >>
rect 96 249 129 257
rect 96 232 104 249
rect 121 232 129 249
rect 96 224 129 232
rect 276 249 309 257
rect 276 232 284 249
rect 301 232 309 249
rect 276 224 309 232
rect 688 249 721 257
rect 688 232 696 249
rect 713 232 721 249
rect 688 224 721 232
rect 801 249 834 257
rect 801 232 809 249
rect 826 232 834 249
rect 801 224 834 232
rect 898 249 931 257
rect 898 232 906 249
rect 923 232 931 249
rect 898 224 931 232
rect 1184 249 1217 257
rect 1184 232 1192 249
rect 1209 232 1217 249
rect 1184 224 1217 232
rect 355 181 388 189
rect 10 164 43 172
rect 10 147 18 164
rect 35 147 43 164
rect 10 139 43 147
rect 62 164 95 172
rect 62 147 70 164
rect 87 147 95 164
rect 62 139 95 147
rect 125 164 158 172
rect 125 147 133 164
rect 150 147 158 164
rect 125 139 158 147
rect 177 164 210 172
rect 177 147 185 164
rect 202 147 210 164
rect 177 139 210 147
rect 240 164 273 172
rect 240 147 248 164
rect 265 147 273 164
rect 240 139 273 147
rect 292 164 325 172
rect 292 147 300 164
rect 317 147 325 164
rect 355 164 363 181
rect 380 164 388 181
rect 355 156 388 164
rect 407 181 440 189
rect 407 164 415 181
rect 432 164 440 181
rect 407 156 440 164
rect 470 181 503 189
rect 470 164 478 181
rect 495 164 503 181
rect 470 156 503 164
rect 522 183 555 189
rect 522 181 615 183
rect 522 164 530 181
rect 547 165 615 181
rect 547 164 555 165
rect 522 156 555 164
rect 292 139 325 147
rect -111 100 -78 108
rect -111 83 -103 100
rect -86 83 -78 100
rect -111 75 -78 83
rect 62 97 82 139
rect 103 98 136 106
rect 103 97 111 98
rect 62 81 111 97
rect 128 81 136 98
rect 305 95 325 139
rect 372 100 405 108
rect 372 95 380 100
rect 62 80 136 81
rect 62 55 82 80
rect 103 73 136 80
rect 184 83 380 95
rect 397 83 405 100
rect 184 75 405 83
rect 184 55 203 75
rect 305 55 325 75
rect 423 55 440 156
rect 496 99 529 107
rect 496 82 504 99
rect 521 82 529 99
rect 496 74 529 82
rect 10 47 43 55
rect 10 30 18 47
rect 35 30 43 47
rect 10 22 43 30
rect 62 47 95 55
rect 62 30 70 47
rect 87 30 95 47
rect 62 22 95 30
rect 125 47 158 55
rect 125 30 133 47
rect 150 30 158 47
rect 125 22 158 30
rect 177 47 210 55
rect 177 30 185 47
rect 202 30 210 47
rect 177 22 210 30
rect 240 47 273 55
rect 240 30 248 47
rect 265 30 273 47
rect 240 22 273 30
rect 292 47 325 55
rect 292 30 300 47
rect 317 30 325 47
rect 292 22 325 30
rect 355 47 388 55
rect 355 30 363 47
rect 380 30 388 47
rect 355 22 388 30
rect 407 50 440 55
rect 407 47 565 50
rect 407 30 415 47
rect 432 30 565 47
rect 407 22 440 30
rect 97 -25 130 -17
rect 97 -42 105 -25
rect 122 -42 130 -25
rect 97 -50 130 -42
rect 214 -25 247 -17
rect 214 -42 222 -25
rect 239 -42 247 -25
rect 214 -50 247 -42
rect 490 -25 523 -17
rect 490 -42 498 -25
rect 515 -42 523 -25
rect 490 -50 523 -42
rect 97 -112 130 -104
rect 97 -129 105 -112
rect 122 -129 130 -112
rect 97 -137 130 -129
rect 210 -112 243 -104
rect 210 -129 218 -112
rect 235 -129 243 -112
rect 210 -137 243 -129
rect 545 -176 565 30
rect 545 -182 574 -176
rect 10 -196 43 -188
rect 10 -213 18 -196
rect 35 -213 43 -196
rect 10 -221 43 -213
rect 62 -196 95 -188
rect 62 -213 70 -196
rect 87 -213 95 -196
rect 62 -221 95 -213
rect 125 -196 158 -188
rect 125 -213 133 -196
rect 150 -213 158 -196
rect 125 -221 158 -213
rect 177 -195 210 -188
rect 240 -195 273 -188
rect 177 -196 273 -195
rect 177 -213 185 -196
rect 202 -213 248 -196
rect 265 -213 273 -196
rect 177 -215 273 -213
rect 177 -221 210 -215
rect 240 -221 273 -215
rect 292 -196 325 -188
rect 292 -213 300 -196
rect 317 -213 325 -196
rect 545 -200 551 -182
rect 568 -200 574 -182
rect 545 -206 574 -200
rect 292 -221 325 -213
rect 65 -270 85 -221
rect 257 -254 290 -246
rect 127 -270 160 -266
rect 65 -274 160 -270
rect 65 -290 135 -274
rect 65 -346 85 -290
rect 127 -291 135 -290
rect 152 -291 160 -274
rect 257 -271 265 -254
rect 282 -271 290 -254
rect 257 -279 290 -271
rect 127 -299 160 -291
rect 308 -300 325 -221
rect 595 -235 615 165
rect 652 164 685 172
rect 652 147 660 164
rect 677 147 685 164
rect 652 139 685 147
rect 704 164 737 172
rect 704 147 712 164
rect 729 147 737 164
rect 704 139 737 147
rect 765 164 798 172
rect 765 147 773 164
rect 790 147 798 164
rect 765 139 798 147
rect 817 164 850 172
rect 817 147 825 164
rect 842 147 850 164
rect 817 139 850 147
rect 717 115 737 139
rect 717 107 800 115
rect 717 95 775 107
rect 654 77 687 85
rect 654 60 662 77
rect 679 60 687 77
rect 654 52 687 60
rect 717 34 737 95
rect 767 90 775 95
rect 792 90 800 107
rect 767 82 800 90
rect 830 83 850 139
rect 923 164 956 172
rect 923 147 931 164
rect 948 147 956 164
rect 923 139 956 147
rect 975 164 1008 172
rect 975 147 983 164
rect 1000 147 1008 164
rect 975 139 1008 147
rect 1036 164 1069 172
rect 1036 147 1044 164
rect 1061 147 1069 164
rect 1036 139 1069 147
rect 1088 164 1121 172
rect 1088 147 1096 164
rect 1113 147 1121 164
rect 1088 139 1121 147
rect 923 100 940 139
rect 988 131 1008 139
rect 958 100 991 105
rect 923 97 991 100
rect 830 77 873 83
rect 830 59 850 77
rect 867 59 873 77
rect 830 53 873 59
rect 923 80 966 97
rect 983 80 991 97
rect 830 35 850 53
rect 652 26 685 34
rect 652 9 660 26
rect 677 9 685 26
rect 652 1 685 9
rect 704 26 737 34
rect 704 9 712 26
rect 729 9 737 26
rect 704 1 737 9
rect 765 27 798 35
rect 765 10 773 27
rect 790 10 798 27
rect 765 2 798 10
rect 817 27 850 35
rect 817 10 825 27
rect 842 10 850 27
rect 817 2 850 10
rect 710 -228 728 1
rect 825 -175 845 2
rect 923 -151 940 80
rect 958 72 991 80
rect 1101 88 1121 139
rect 1195 163 1228 171
rect 1195 146 1203 163
rect 1220 146 1228 163
rect 1195 138 1228 146
rect 1247 163 1280 171
rect 1247 146 1255 163
rect 1272 146 1280 163
rect 1247 138 1280 146
rect 1144 95 1177 103
rect 1144 88 1152 95
rect 1101 78 1152 88
rect 1169 78 1177 95
rect 1101 70 1177 78
rect 1032 56 1065 64
rect 1032 39 1040 56
rect 1057 39 1065 56
rect 1032 31 1065 39
rect 1065 -51 1085 -44
rect 1005 -59 1038 -51
rect 1005 -76 1013 -59
rect 1030 -76 1038 -59
rect 1005 -84 1038 -76
rect 1057 -59 1090 -51
rect 1157 -55 1177 70
rect 1247 96 1267 138
rect 1294 97 1323 103
rect 1294 96 1300 97
rect 1247 79 1300 96
rect 1317 79 1323 97
rect 1247 54 1267 79
rect 1294 73 1323 79
rect 1195 46 1228 54
rect 1195 29 1203 46
rect 1220 29 1228 46
rect 1195 21 1228 29
rect 1247 46 1280 54
rect 1247 29 1255 46
rect 1272 29 1280 46
rect 1247 21 1280 29
rect 1275 -23 1308 -15
rect 1275 -40 1283 -23
rect 1300 -40 1308 -23
rect 1275 -48 1308 -40
rect 1057 -76 1065 -59
rect 1082 -76 1090 -59
rect 1057 -84 1090 -76
rect 1117 -77 1177 -55
rect 977 -151 997 -144
rect 1060 -150 1079 -84
rect 1117 -150 1137 -77
rect 917 -159 950 -151
rect 765 -183 798 -175
rect 765 -200 773 -183
rect 790 -200 798 -183
rect 765 -208 798 -200
rect 817 -183 850 -175
rect 817 -200 825 -183
rect 842 -200 850 -183
rect 917 -176 925 -159
rect 942 -176 950 -159
rect 917 -184 950 -176
rect 969 -155 1002 -151
rect 1057 -155 1090 -150
rect 969 -158 1090 -155
rect 969 -159 1065 -158
rect 969 -176 977 -159
rect 994 -175 1065 -159
rect 1082 -175 1090 -158
rect 994 -176 1002 -175
rect 969 -184 1002 -176
rect 1057 -183 1090 -175
rect 1109 -158 1142 -150
rect 1109 -175 1117 -158
rect 1134 -175 1142 -158
rect 1109 -183 1142 -175
rect 1065 -185 1085 -183
rect 817 -208 850 -200
rect 1083 -212 1116 -204
rect 943 -221 976 -213
rect 651 -235 684 -228
rect 423 -236 684 -235
rect 423 -253 659 -236
rect 676 -253 684 -236
rect 423 -255 684 -253
rect 372 -299 405 -291
rect 372 -300 380 -299
rect 185 -316 380 -300
rect 397 -316 405 -299
rect 185 -320 405 -316
rect 185 -346 205 -320
rect 245 -346 265 -339
rect 302 -346 320 -320
rect 372 -324 405 -320
rect 423 -346 440 -255
rect 651 -261 684 -255
rect 703 -236 736 -228
rect 703 -253 711 -236
rect 728 -253 736 -236
rect 943 -238 951 -221
rect 968 -238 976 -221
rect 1083 -229 1091 -212
rect 1108 -229 1116 -212
rect 1083 -237 1116 -229
rect 943 -246 976 -238
rect 703 -261 736 -253
rect 660 -322 678 -261
rect 790 -278 823 -270
rect 790 -295 798 -278
rect 815 -295 823 -278
rect 790 -303 823 -295
rect 1086 -322 1105 -237
rect 660 -341 1105 -322
rect 10 -354 43 -346
rect 10 -371 18 -354
rect 35 -371 43 -354
rect 10 -379 43 -371
rect 62 -354 95 -346
rect 62 -371 70 -354
rect 87 -371 95 -354
rect 62 -379 95 -371
rect 125 -354 158 -346
rect 125 -371 133 -354
rect 150 -371 158 -354
rect 125 -379 158 -371
rect 177 -354 210 -346
rect 177 -371 185 -354
rect 202 -371 210 -354
rect 177 -379 210 -371
rect 240 -354 273 -346
rect 240 -371 248 -354
rect 265 -371 273 -354
rect 240 -379 273 -371
rect 292 -354 325 -346
rect 292 -371 300 -354
rect 317 -371 325 -354
rect 292 -379 325 -371
rect 355 -354 388 -346
rect 355 -371 363 -354
rect 380 -371 388 -354
rect 355 -379 388 -371
rect 407 -354 440 -346
rect 407 -371 415 -354
rect 432 -371 440 -354
rect 407 -379 440 -371
rect 94 -423 127 -415
rect 94 -440 102 -423
rect 119 -440 127 -423
rect 94 -448 127 -440
rect 249 -423 282 -415
rect 249 -440 257 -423
rect 274 -440 282 -423
rect 249 -448 282 -440
<< viali >>
rect 104 232 121 249
rect 284 232 301 249
rect 696 232 713 249
rect 809 232 826 249
rect 906 232 923 249
rect 1192 232 1209 249
rect 18 147 35 164
rect 70 147 87 164
rect 133 147 150 164
rect 185 147 202 164
rect 248 147 265 164
rect 300 147 317 164
rect 363 164 380 181
rect 415 164 432 181
rect 478 164 495 181
rect 530 164 547 181
rect -103 83 -86 100
rect 111 81 128 98
rect 380 83 397 100
rect 504 82 521 99
rect 18 30 35 47
rect 70 30 87 47
rect 133 30 150 47
rect 185 30 202 47
rect 248 30 265 47
rect 300 30 317 47
rect 363 30 380 47
rect 415 30 432 47
rect 105 -42 122 -25
rect 222 -42 239 -25
rect 498 -42 515 -25
rect 105 -129 122 -112
rect 218 -129 235 -112
rect 18 -213 35 -196
rect 70 -213 87 -196
rect 133 -213 150 -196
rect 185 -213 202 -196
rect 248 -213 265 -196
rect 300 -213 317 -196
rect 551 -200 568 -182
rect 135 -291 152 -274
rect 265 -271 282 -254
rect 660 147 677 164
rect 712 147 729 164
rect 773 147 790 164
rect 825 147 842 164
rect 662 60 679 77
rect 931 147 948 164
rect 983 147 1000 164
rect 1044 147 1061 164
rect 1096 147 1113 164
rect 850 59 867 77
rect 966 80 983 97
rect 660 9 677 26
rect 712 9 729 26
rect 773 10 790 27
rect 825 10 842 27
rect 1203 146 1220 163
rect 1255 146 1272 163
rect 1152 78 1169 95
rect 1040 39 1057 56
rect 1013 -76 1030 -59
rect 1300 79 1317 97
rect 1203 29 1220 46
rect 1255 29 1272 46
rect 1283 -40 1300 -23
rect 1065 -76 1082 -59
rect 773 -200 790 -183
rect 825 -200 842 -183
rect 925 -176 942 -159
rect 977 -176 994 -159
rect 1065 -175 1082 -158
rect 1117 -175 1134 -158
rect 659 -253 676 -236
rect 380 -316 397 -299
rect 711 -253 728 -236
rect 951 -238 968 -221
rect 1091 -229 1108 -212
rect 798 -295 815 -278
rect 18 -371 35 -354
rect 70 -371 87 -354
rect 133 -371 150 -354
rect 185 -371 202 -354
rect 248 -371 265 -354
rect 300 -371 317 -354
rect 363 -371 380 -354
rect 415 -371 432 -354
rect 102 -440 119 -423
rect 257 -440 274 -423
<< metal1 >>
rect -10 250 948 257
rect -48 249 948 250
rect -48 232 104 249
rect 121 232 284 249
rect 301 232 696 249
rect 713 232 809 249
rect 826 232 906 249
rect 923 242 948 249
rect 1174 249 1227 257
rect 1174 242 1192 249
rect 923 232 1192 242
rect 1209 232 1227 249
rect -48 231 1227 232
rect -111 100 -78 108
rect -111 83 -103 100
rect -86 83 -78 100
rect -111 75 -78 83
rect -48 -104 -25 231
rect -10 224 1227 231
rect 20 172 40 224
rect 135 172 155 224
rect 365 189 385 224
rect 475 189 495 224
rect 355 181 388 189
rect 10 164 43 172
rect 10 147 18 164
rect 35 147 43 164
rect 10 139 43 147
rect 62 164 95 172
rect 62 147 70 164
rect 87 147 95 164
rect 62 139 95 147
rect 125 164 158 172
rect 125 147 133 164
rect 150 147 158 164
rect 125 139 158 147
rect 177 170 210 172
rect 240 170 273 172
rect 177 164 273 170
rect 177 147 185 164
rect 202 150 248 164
rect 202 147 210 150
rect 177 139 210 147
rect 240 147 248 150
rect 265 147 273 164
rect 240 139 273 147
rect 292 164 325 172
rect 292 147 300 164
rect 317 147 325 164
rect 355 164 363 181
rect 380 164 388 181
rect 355 156 388 164
rect 407 181 440 189
rect 407 164 415 181
rect 432 164 440 181
rect 407 156 440 164
rect 470 181 503 189
rect 470 164 478 181
rect 495 164 503 181
rect 470 156 503 164
rect 522 181 555 189
rect 522 164 530 181
rect 547 164 555 181
rect 655 172 675 224
rect 765 172 785 224
rect 926 172 946 186
rect 1036 172 1056 224
rect 1205 185 1224 224
rect 522 156 555 164
rect 652 164 685 172
rect 292 139 325 147
rect 652 147 660 164
rect 677 147 685 164
rect 652 139 685 147
rect 704 164 737 172
rect 704 147 712 164
rect 729 147 737 164
rect 704 139 737 147
rect 765 164 798 172
rect 765 147 773 164
rect 790 147 798 164
rect 765 139 798 147
rect 817 164 850 172
rect 817 147 825 164
rect 842 147 850 164
rect 817 139 850 147
rect 923 164 956 172
rect 923 147 931 164
rect 948 147 956 164
rect 923 139 956 147
rect 975 164 1008 172
rect 975 147 983 164
rect 1000 147 1008 164
rect 975 139 1008 147
rect 1036 164 1069 172
rect 1036 147 1044 164
rect 1061 147 1069 164
rect 1036 139 1069 147
rect 1088 164 1121 172
rect 1205 171 1225 185
rect 1088 147 1096 164
rect 1113 147 1121 164
rect 1088 139 1121 147
rect 1195 163 1228 171
rect 1195 146 1203 163
rect 1220 146 1228 163
rect 1195 138 1228 146
rect 1247 163 1280 171
rect 1247 146 1255 163
rect 1272 146 1280 163
rect 1247 138 1280 146
rect 103 98 136 106
rect 103 81 111 98
rect 128 81 136 98
rect 103 73 136 81
rect 372 100 405 108
rect 372 83 380 100
rect 397 83 405 100
rect 372 75 405 83
rect 496 99 529 107
rect 496 82 504 99
rect 521 82 529 99
rect 958 97 991 105
rect 496 74 529 82
rect 654 77 687 85
rect 10 47 43 55
rect 10 30 18 47
rect 35 30 43 47
rect 10 22 43 30
rect 62 47 95 55
rect 62 30 70 47
rect 87 30 95 47
rect 62 22 95 30
rect 125 47 158 55
rect 125 30 133 47
rect 150 30 158 47
rect 125 22 158 30
rect 177 47 210 55
rect 177 30 185 47
rect 202 30 210 47
rect 177 22 210 30
rect 240 47 273 55
rect 240 30 248 47
rect 265 30 273 47
rect 240 22 273 30
rect 292 47 325 55
rect 292 30 300 47
rect 317 30 325 47
rect 292 22 325 30
rect 355 47 388 55
rect 355 30 363 47
rect 380 30 388 47
rect 355 22 388 30
rect 407 47 440 55
rect 407 30 415 47
rect 432 30 440 47
rect 407 22 440 30
rect 23 -17 43 22
rect 135 -17 155 22
rect 248 -17 268 22
rect 300 20 320 22
rect 360 -17 380 22
rect 501 -16 520 74
rect 654 60 662 77
rect 679 75 687 77
rect 844 77 873 83
rect 844 75 850 77
rect 679 60 850 75
rect 654 59 850 60
rect 867 59 873 77
rect 958 80 966 97
rect 983 80 991 97
rect 958 72 991 80
rect 1144 95 1177 103
rect 1144 78 1152 95
rect 1169 78 1177 95
rect 1144 70 1177 78
rect 1294 97 1323 103
rect 1294 79 1300 97
rect 1317 79 1323 97
rect 1294 73 1323 79
rect 654 55 873 59
rect 654 52 687 55
rect 844 53 873 55
rect 1032 56 1065 64
rect 1032 39 1040 56
rect 1057 39 1065 56
rect 652 26 685 34
rect 652 9 660 26
rect 677 9 685 26
rect 652 1 685 9
rect 704 26 737 34
rect 704 9 712 26
rect 729 9 737 26
rect 704 1 737 9
rect 765 27 798 35
rect 765 10 773 27
rect 790 10 798 27
rect 765 2 798 10
rect 817 27 850 35
rect 1032 31 1065 39
rect 1195 46 1228 54
rect 817 10 825 27
rect 842 10 850 27
rect 1195 29 1203 46
rect 1220 29 1228 46
rect 1195 21 1228 29
rect 1247 46 1280 54
rect 1247 29 1255 46
rect 1272 29 1280 46
rect 1247 21 1280 29
rect 817 2 850 10
rect 1200 19 1228 21
rect 655 -1 677 1
rect 655 -16 675 -1
rect 770 -16 790 2
rect 1200 -15 1219 19
rect 886 -16 1312 -15
rect 501 -17 1312 -16
rect 15 -23 1312 -17
rect 15 -25 1283 -23
rect 15 -42 105 -25
rect 122 -42 222 -25
rect 239 -42 498 -25
rect 515 -35 1283 -25
rect 515 -42 1030 -35
rect 15 -50 1030 -42
rect 1271 -40 1283 -35
rect 1300 -40 1312 -23
rect 1271 -48 1312 -40
rect -48 -112 350 -104
rect -48 -129 105 -112
rect 122 -129 218 -112
rect 235 -129 350 -112
rect -48 -137 350 -129
rect 15 -188 35 -137
rect 135 -188 155 -137
rect 10 -196 43 -188
rect 10 -213 18 -196
rect 35 -213 43 -196
rect 10 -221 43 -213
rect 62 -196 95 -188
rect 62 -213 70 -196
rect 87 -213 95 -196
rect 62 -221 95 -213
rect 125 -196 158 -188
rect 125 -213 133 -196
rect 150 -213 158 -196
rect 125 -221 158 -213
rect 177 -196 210 -188
rect 177 -213 185 -196
rect 202 -213 210 -196
rect 177 -221 210 -213
rect 240 -196 273 -188
rect 240 -213 248 -196
rect 265 -213 273 -196
rect 240 -221 273 -213
rect 292 -196 325 -188
rect 292 -213 300 -196
rect 317 -213 325 -196
rect 292 -221 325 -213
rect 257 -254 290 -246
rect 127 -274 160 -266
rect 127 -291 135 -274
rect 152 -291 160 -274
rect 257 -271 265 -254
rect 282 -271 290 -254
rect 257 -279 290 -271
rect 127 -299 160 -291
rect 372 -299 405 -291
rect 372 -316 380 -299
rect 397 -316 405 -299
rect 372 -324 405 -316
rect 10 -354 43 -346
rect 10 -371 18 -354
rect 35 -371 43 -354
rect 10 -379 43 -371
rect 62 -354 95 -346
rect 62 -371 70 -354
rect 87 -371 95 -354
rect 62 -379 95 -371
rect 125 -354 158 -346
rect 125 -371 133 -354
rect 150 -371 158 -354
rect 125 -379 158 -371
rect 177 -354 210 -346
rect 177 -371 185 -354
rect 202 -371 210 -354
rect 177 -379 210 -371
rect 240 -354 273 -346
rect 240 -371 248 -354
rect 265 -371 273 -354
rect 240 -379 273 -371
rect 292 -354 325 -346
rect 292 -371 300 -354
rect 317 -371 325 -354
rect 292 -379 325 -371
rect 355 -354 388 -346
rect 355 -371 363 -354
rect 380 -371 388 -354
rect 355 -379 388 -371
rect 407 -354 440 -346
rect 407 -371 415 -354
rect 432 -371 440 -354
rect 407 -379 440 -371
rect 15 -415 35 -379
rect 140 -415 158 -379
rect 248 -415 268 -379
rect 300 -381 320 -379
rect 365 -415 385 -379
rect 456 -415 475 -50
rect 1005 -51 1030 -50
rect 1005 -59 1038 -51
rect 1005 -76 1013 -59
rect 1030 -76 1038 -59
rect 1005 -84 1038 -76
rect 1057 -59 1090 -51
rect 1057 -76 1065 -59
rect 1082 -76 1090 -59
rect 1057 -84 1090 -76
rect 1010 -86 1030 -84
rect 917 -159 950 -151
rect 545 -182 574 -176
rect 545 -200 551 -182
rect 568 -185 574 -182
rect 765 -183 798 -175
rect 765 -185 773 -183
rect 568 -200 773 -185
rect 790 -200 798 -183
rect 545 -205 798 -200
rect 545 -206 574 -205
rect 765 -208 798 -205
rect 817 -183 850 -175
rect 817 -200 825 -183
rect 842 -200 850 -183
rect 917 -176 925 -159
rect 942 -176 950 -159
rect 917 -184 950 -176
rect 969 -159 1002 -151
rect 969 -176 977 -159
rect 994 -176 1002 -159
rect 969 -184 1002 -176
rect 1057 -158 1090 -150
rect 1057 -175 1065 -158
rect 1082 -175 1090 -158
rect 1057 -183 1090 -175
rect 1109 -158 1142 -150
rect 1109 -175 1117 -158
rect 1134 -175 1142 -158
rect 1109 -183 1142 -175
rect 922 -186 942 -184
rect 1062 -185 1082 -183
rect 817 -208 850 -200
rect 770 -210 790 -208
rect 770 -227 789 -210
rect 1083 -212 1116 -204
rect 943 -221 976 -213
rect 943 -227 951 -221
rect 651 -236 684 -228
rect 651 -253 659 -236
rect 676 -253 684 -236
rect 651 -261 684 -253
rect 703 -236 736 -228
rect 703 -253 711 -236
rect 728 -253 736 -236
rect 770 -238 951 -227
rect 968 -238 976 -221
rect 1083 -229 1091 -212
rect 1108 -229 1116 -212
rect 1083 -237 1116 -229
rect 770 -246 976 -238
rect 703 -261 736 -253
rect 656 -263 676 -261
rect 790 -278 823 -270
rect 790 -295 798 -278
rect 815 -295 823 -278
rect 790 -303 823 -295
rect -52 -423 475 -415
rect -52 -440 102 -423
rect 119 -440 257 -423
rect 274 -440 475 -423
rect -52 -448 475 -440
<< labels >>
flabel locali s -98 87 -90 96 0 FreeSans 400 0 0 0 din
port 0 nsew
flabel locali s 269 -268 277 -259 0 FreeSans 400 0 0 0 wb
port 1 nsew
flabel metal1 s 107 -436 115 -427 0 FreeSans 400 0 0 0 gnd
port 2 nsew
flabel metal1 s 108 237 116 246 0 FreeSans 400 0 0 0 vdd
port 3 nsew
flabel locali s 420 36 428 45 0 FreeSans 400 0 0 0 blb
port 4 nsew
flabel locali s 536 168 544 177 0 FreeSans 400 0 0 0 bl
port 5 nsew
flabel locali s 666 64 674 73 0 FreeSans 400 0 0 0 qb
port 6 nsew
flabel locali s 779 95 787 104 0 FreeSans 400 0 0 0 q
port 7 nsew
flabel locali s 800 -292 808 -283 0 FreeSans 400 0 0 0 wl
port 8 nsew
flabel locali s 1045 42 1053 51 0 FreeSans 400 0 0 0 rd_en
port 9 nsew
flabel locali s 1302 85 1310 94 0 FreeSans 400 0 0 0 dout
port 10 nsew
flabel locali 72 84 79 92 0 FreeSans 200 0 0 0 net1
flabel locali 310 81 317 89 0 FreeSans 200 0 0 0 net2
flabel metal1 218 157 225 165 0 FreeSans 200 0 0 0 net3
flabel locali 71 -285 78 -277 0 FreeSans 200 0 0 0 net4
flabel locali 308 -312 315 -304 0 FreeSans 200 0 0 0 net5
flabel locali 930 83 947 91 0 FreeSans 200 0 0 0 net6
flabel locali 1106 74 1123 82 0 FreeSans 200 0 0 0 net7
flabel locali 1068 -124 1075 -105 0 FreeSans 200 0 0 0 net8
flabel locali 217 -210 231 -204 0 FreeSans 200 0 0 0 net9
<< end >>
